module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input LIOB33_X0Y123_IOB_X0Y124_IPAD,
  input LIOB33_X0Y125_IOB_X0Y125_IPAD,
  input LIOB33_X0Y125_IOB_X0Y126_IPAD,
  input LIOB33_X0Y127_IOB_X0Y127_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CMUX;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AMUX;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_DO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_CO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_DO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AMUX;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_AMUX;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_AO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_BO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_BO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_CO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_CO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_DO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_DO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e800ff008000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f88880000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000120002000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fecc0000cccc)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_BLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h050505050000a000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee888888880000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcffffffff)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc550000cc550c05)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I5(LIOB33_X0Y123_IOB_X0Y123_I),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000100)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_DO6),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f0101011111111)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33000000ff000f00)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y121_IOB_X0Y121_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000b0300000f0f)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(LIOB33_X0Y127_IOB_X0Y127_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h40c040c0440050f0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y127_IOB_X0Y127_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h220000000a000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffaaafaaaf)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_DO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffffffffffff)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_BLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0fcfffff5fd)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_CO6),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_BO6),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30300000f0ff0000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(LIOB33_X0Y121_IOB_X0Y121_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_DO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_CO6),
.I3(CLBLL_L_X2Y116_SLICE_X0Y116_BO6),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffcdffffffff)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I5(CLBLL_L_X2Y116_SLICE_X0Y116_BO6),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001010100)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_ALUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_DO6),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(CLBLL_L_X2Y116_SLICE_X0Y116_CO6),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff00000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(1'b1),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(LIOB33_X0Y121_IOB_X0Y122_I),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0e0c0e0c)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_BO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000f000e0)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800080000008800)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffa0a0a0a0)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3322332333333333)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_BO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff04ffaaffaeff)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeeeeeeeeeeee)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(RIOB33_X105Y119_IOB_X1Y120_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h01cd00000dcd0000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050004)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_DO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fffffffff7ffff)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f11111f5f1111)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_DO6),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeeeeeeeaee)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y119_IOB_X0Y120_I),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfff0b3b3b3b3)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y127_IOB_X0Y127_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef8f8f000000011)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555455555)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I1(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(LIOB33_X0Y125_IOB_X0Y125_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ea00c000ff00ff)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300220003000200)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80800000ff80ff00)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y119_IOB_X1Y120_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X2Y114_SLICE_X1Y114_CO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222222ff22ff)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f4005400000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff88ffaaffa8)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I3(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafa00a0000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(1'b1),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_DO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_CO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_BO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_DO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_CO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_BO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffbbffbfffffff)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_ALUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_DO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_CO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_BO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4f4f455555555)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_ALUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_AO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_DO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_CO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_BO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_AO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000088000000ff)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(1'b1),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33fb33fb00fa00fa)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff0001)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff5dffff)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f4ffffffff)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000010000ffbb)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5010551100000000)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfffffffdfd)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaeeeeeeeeeeeec)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000aa20)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0707070f88888800)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000302000002000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y127_IOB_X0Y127_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000013)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I4(CLBLL_L_X2Y116_SLICE_X1Y116_BO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc00fcfcfc00fc54)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.I2(LIOB33_X0Y127_IOB_X0Y127_I),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha800fcfcfcfcfcfc)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfccccffdffcdc)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y124_I),
.I1(LIOB33_X0Y123_IOB_X0Y123_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f0fff03322ff22)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000fffff000f222f)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff444444ff4cfcfc)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(LIOB33_X0Y127_IOB_X0Y127_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f000bbbbabbb)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500550055)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h008cdc8c00040404)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y125_IOB_X0Y125_I),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d5d5c000d555)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff11f111f1)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.I1(RIOB33_X105Y119_IOB_X1Y120_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff030ffffa020)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.I1(RIOB33_X105Y119_IOB_X1Y120_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.I5(RIOB33_X105Y119_IOB_X1Y119_I),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbafbf00000000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3fffffcfcacf0a)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa0000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333330030303000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.I5(LIOB33_X0Y125_IOB_X0Y125_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777707077007000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000feeefaaa)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_BO6),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0e000000011)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccefccefcc)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLL_L_X2Y113_SLICE_X1Y113_CO6),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005500ff0f5505)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(1'b1),
.I2(LIOB33_X0Y127_IOB_X0Y127_I),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7f3f3f77ff33ff)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb00bb0000000b00)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0fdfcf5500ddcc)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffbfffffffb)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222fff2ffffffff)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffddfffcff)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00010001fffe0000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f7f0f077f700f0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0002000a000a00)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I1(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0700000000000000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a3000300030003)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y124_I),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(LIOB33_X0Y121_IOB_X0Y122_I),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f3f7f3f5f0f5f0f)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffffefeffff)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLL_L_X2Y114_SLICE_X1Y114_BO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfdddfdddddddff)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00feaaaafefe)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h08000a0008080a0a)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3000301000000010)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77f070fffff0f0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff01ff00000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3b0a3b3b)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00880000008a0000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_AO6),
.I5(LIOB33_X0Y121_IOB_X0Y122_I),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccccffdcff)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_CO6),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y121_IOB_X0Y121_I),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0d0d0d000dd00dd)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(LIOB33_X0Y123_IOB_X0Y124_I),
.I1(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0ffeefffe)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(LIOB33_X0Y127_IOB_X0Y127_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y123_IOB_X0Y123_I),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fff077005550)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3322333303020303)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y127_IOB_X0Y127_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1110000011101110)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100cdcc0300cfcc)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcffffa8fca8fc)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0c3f3f00000030)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(1'b1),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffccffffffff)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff4044444040)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y121_IOB_X0Y121_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000110000cfcccf)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444440000cc0088)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(1'b1),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h003f00ffffffffff)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfefe00cc00fe)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555500ffdfdfcfff)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0000044404400)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLL_L_X2Y116_SLICE_X1Y116_BO6),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000b0b1bbbb)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I2(CLBLL_L_X2Y119_SLICE_X1Y119_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000332200000302)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000d5d5d5dd)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e0e0e0c0c0c0c)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffee55545544)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f1f5f0f5f0f5f0)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_DO6),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff32ffffff33ffff)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0eeeeee00eeeeee)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f7fffffdfff5f5f)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5755ffff5555)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff8850)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h004400440000f2f0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000100000000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.I2(CLBLL_L_X2Y116_SLICE_X1Y116_BO6),
.I3(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.I4(1'b1),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005000400000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I1(CLBLL_L_X2Y116_SLICE_X1Y116_CO6),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f0f5f1f1f5f5)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f5f5000000ff)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccfffafac8fa)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000002)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3330fffc3330fffd)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000af0000008c)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0055ffff0050)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a00000002)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0a3f3b0f0a0f0a)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_CO6),
.I1(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00af00ccffdcff)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff57575757)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555111155441100)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333000033320000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0100000101)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5655000055550000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000abaaaaaa)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000ff00ff)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555554455ff5555)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000a08)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff33333332)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0b0f0f0f0a)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00dc8c8c00040404)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y124_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y126_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y127_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y116_SLICE_X0Y116_DO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X1Y117_DO6),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_DO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X2Y143_SLICE_X0Y143_AO5),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X2Y129_SLICE_X0Y129_AO5),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLL_L_X2Y143_SLICE_X0Y143_AO6),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_AMUX = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_BMUX = CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_AMUX = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_AMUX = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_AMUX = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_BMUX = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_CMUX = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D = CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_AMUX = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_AMUX = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_AMUX = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_AMUX = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_AMUX = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_BMUX = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AMUX = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_AMUX = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B = CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D = CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B = CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C = CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D = CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B = CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D = CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_AMUX = CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A = CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B = CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D = CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A = CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B = CLBLL_L_X2Y143_SLICE_X0Y143_BO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C = CLBLL_L_X2Y143_SLICE_X0Y143_CO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D = CLBLL_L_X2Y143_SLICE_X0Y143_DO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_AMUX = CLBLL_L_X2Y143_SLICE_X0Y143_AO5;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A = CLBLL_L_X2Y143_SLICE_X1Y143_AO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B = CLBLL_L_X2Y143_SLICE_X1Y143_BO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C = CLBLL_L_X2Y143_SLICE_X1Y143_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D = CLBLL_L_X2Y143_SLICE_X1Y143_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AMUX = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_AMUX = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_AMUX = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_AMUX = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_BMUX = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AMUX = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_AMUX = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AMUX = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_AMUX = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CMUX = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AMUX = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_AMUX = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_AMUX = CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_BMUX = CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_AMUX = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_CMUX = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_DMUX = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_AMUX = CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_BMUX = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_AMUX = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_AMUX = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_BMUX = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_AMUX = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_BMUX = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_AMUX = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_AMUX = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_BMUX = CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_AMUX = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X2Y143_SLICE_X0Y143_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A5 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A6 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B5 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A4 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A1 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A4 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A2 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A3 = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A4 = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A5 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A6 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D5 = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D6 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A1 = CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A3 = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A4 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B1 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B5 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B6 = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C2 = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C3 = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C4 = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C5 = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D4 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X2Y143_SLICE_X0Y143_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A1 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A3 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B6 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C6 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D6 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A3 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A5 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X2Y143_SLICE_X0Y143_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
endmodule
