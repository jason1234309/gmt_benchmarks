module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AMUX;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AMUX;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BMUX;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_AMUX;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_AO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_BMUX;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_BO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_CO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_CO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_DO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_DO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_BO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_BO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_DO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_DO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AMUX;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AMUX;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CMUX;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CLK;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B5Q;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CLK;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A5Q;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5Q;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5Q;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B5Q;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B5Q;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CLK;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CLK;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CLK;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CLK;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DMUX;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CLK;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AMUX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BMUX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C5Q;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CLK;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CMUX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_DO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CLK;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A5Q;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AMUX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CLK;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_DO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CLK;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B5Q;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BMUX;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C5Q;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CLK;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CMUX;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A5Q;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AMUX;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B5Q;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BMUX;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CLK;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A5Q;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CLK;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CLK;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CLK;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CLK;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A5Q;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AMUX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CLK;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CMUX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CLK;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DMUX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CLK;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CLK;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CE;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CLK;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_SR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CLK;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D5Q;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CLK;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CLK;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B5Q;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CLK;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CLK;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CE;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CLK;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_SR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CE;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CLK;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_SR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CLK;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CMUX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DMUX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CLK;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CMUX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_DO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CLK;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_DO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CLK;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BMUX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CLK;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_DO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_DO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_BO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_BO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_CO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_CO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_DO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_DO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_AO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_BO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_BO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_CO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_CO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_DO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_DO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_AO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_AO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_BO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_BO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_CO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_CO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_DO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_DO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AMUX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_DO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_DO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_AO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_AO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_BO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_BO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_CO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_CO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_DO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_DO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A5Q;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C5Q;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A5Q;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5Q;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5Q;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5Q;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CLK;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CLK;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DMUX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_AO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_AO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_BO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_BO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_CO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_CO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_DO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_DO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AMUX;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_BO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_BO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_CO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_CO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_DO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_DO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AMUX;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AMUX;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CLK;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CLK;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CLK;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CLK;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A5Q;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B5Q;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B5Q;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C5Q;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CLK;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CLK;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CLK;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CLK;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CLK;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CLK;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CLK;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CLK;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D5Q;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A5Q;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CLK;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CLK;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CLK;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BMUX;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CLK;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CLK;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CLK;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_AO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_AO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_BO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_BO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CLK;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_DO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_DO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_BO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_BO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_CO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_CO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_DO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_DO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A5Q;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AMUX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AQ;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BMUX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_CLK;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_DO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_DO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CLK;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_DO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_DO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A5Q;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AMUX;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AQ;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AX;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_BO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_BO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_BQ;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_CLK;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_CO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_CO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_CQ;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_DO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_DO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_AO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_AO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_BO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_BO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_CO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_CO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_DO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_DO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_AO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_BO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_BO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_CLK;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_CO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_DO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_DO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_AO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_AO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_AQ;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_BO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_BO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_BQ;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_CLK;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_CMUX;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_CO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_CO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_DO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_DO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DMUX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_BO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_BO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_CO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_DO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_DO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AQ;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BQ;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CLK;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CQ;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DQ;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_AO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_AO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_AQ;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_BO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_BO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_BQ;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_CLK;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_CO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_CQ;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_DO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AQ;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BMUX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CLK;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CQ;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_DO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_AQ;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_BO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_BO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_CLK;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_CO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_CO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_DO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_DO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AQ;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BQ;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CLK;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CQ;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_DMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_DO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_DO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_AO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_BO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_CO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_DO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_DO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A5Q;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AMUX;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AQ;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AX;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_BO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_BO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_BQ;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CLK;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CQ;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_DMUX;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_DO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_AO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_AO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_AQ;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_AX;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_BO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_CLK;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_CO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_CO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_DO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_DO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CLK;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_DO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_DO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_AMUX;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_AO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_BO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_CO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_CO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_DO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_DO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_BO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_BO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_CO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_CO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_DO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_DO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_AO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_AO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_BO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_BO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CLK;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CQ;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_DO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_AMUX;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_AO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_AO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_BO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_CO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_DO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_DO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_BMUX;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CLK;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_DO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_DO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_AO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_AO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_BO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_BO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_CO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_DO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_DO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_AO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_AO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_AQ;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_BO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_BO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CLK;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_DO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_DO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_AO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_BO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_CO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_DO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_DO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CLK;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_DO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_BO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_CO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_DO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D_XOR;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A1;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A2;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A3;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A4;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_AO5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_AO6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A_CY;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_A_XOR;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B1;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B2;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B3;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B4;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_BO5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_BO6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B_CY;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_B_XOR;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C1;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C2;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C3;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C4;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_CO5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_CO6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C_CY;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_C_XOR;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D1;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D2;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D3;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D4;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_DO5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_DO6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D_CY;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X56Y143_D_XOR;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A1;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A2;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A3;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A4;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_AO5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_AO6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A_CY;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_A_XOR;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B1;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B2;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B3;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B4;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_BO5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_BO6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B_CY;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_B_XOR;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C1;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C2;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C3;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C4;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_CO5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_CO6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C_CY;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_C_XOR;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D1;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D2;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D3;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D4;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_DO5;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_DO6;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D_CY;
  wire [0:0] CLBLM_R_X37Y143_SLICE_X57Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CLK;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BMUX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5Q;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CLK;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CLK;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CLK;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B5Q;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D5Q;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y138_SLICE_X4Y138_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc0f000f00)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I2(CLBLL_L_X4Y138_SLICE_X4Y138_AO6),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfbfffbfffb)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefffffefeffff)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_DO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_CO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefffffffeeffff)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_BO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffffffeeffff)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_AO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_DO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_CO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_BO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_AO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h030b000a030b000a)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_BLUT (
.I0(LIOB33_X0Y55_IOB_X0Y55_I),
.I1(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.I4(LIOB33_X0Y71_IOB_X0Y71_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h030b000a030b000a)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffff33ffffff)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000400040f0f0004)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_ALUT (
.I0(CLBLL_L_X2Y147_SLICE_X0Y147_AO5),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_B5Q),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbfffff)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0001010101)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbffffbffff)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88ff8888f8fff8f8)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.I1(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff80000ff880000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I2(LIOB33_X0Y53_IOB_X0Y53_I),
.I3(CLBLL_L_X4Y138_SLICE_X4Y138_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_DO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_AO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_CO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888d8800005500)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabeaa00001400)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_AO5),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_A5Q),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3a0eca0eca0eca0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_DO5),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcddc0110cccc0000)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_AO6),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880088008800)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_BLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800080000000)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_DO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_AO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_BO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_CO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf088880000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_AO5),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habaa0100aeaa0400)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.I2(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00006ccc6ccc)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff48c048c048c0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_DO5),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_AO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_BO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf070f03055550000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_CLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_D5Q),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.I4(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfafa0a0a)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_BLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.I1(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I5(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33333030)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_ALUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_AO6),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011000000130000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_CO6),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001414ff000000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_BO6),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_CO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f5f7f7f5f5f5f5)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_D5Q),
.I4(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aca0a3a0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_CLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00c3aaaa0000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_BLUT (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_AO6),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff5a005a)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444cccc5555ffff)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_BQ),
.I1(CLBLM_R_X13Y142_SLICE_X18Y142_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00007f7f7f7f)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_DO6),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffffffffffff)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_BLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_CO6),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fff0fffdfff5fff)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_ALUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_DO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf05acccc0000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y141_SLICE_X4Y141_CO6),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f088880000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_CLUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.I2(RIOB33_X105Y127_IOB_X1Y127_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f03300cc00)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14fa50aa00aa00)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbbffbbff)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_CO6),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00000000000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_CO6),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hba30ba30bb33ba30)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_ALUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I3(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_DQ),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0cc0aaaa0cc0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_AO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_BO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05550fffffffffff)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_DLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff135f80008000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_CLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_DQ),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfc0cfc0c0c0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aaffaa30aaf0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_ALUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_AO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_BO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000054045404)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffffffdf)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00fff0f0aaaa)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_BQ),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff28a0000028a0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_DQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X5Y145_AO6),
.Q(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044554400)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b3bff3b0a0aff0a)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_CLUT (
.I0(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h73ff737350ff5050)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.I2(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.I4(CLBLM_L_X12Y141_SLICE_X16Y141_C5Q),
.I5(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f3f3ff00c0c0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I2(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff22fff2)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_DLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.I2(LIOB33_X0Y65_IOB_X0Y65_I),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_AO5),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_DO6),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffddfdccfc)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.I5(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3f3a2a2a2a2)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_ALUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_B5Q),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(1'b1),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00afaaafaa)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_DLUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff2f2f2222)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.I5(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccfceefe)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_AO6),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_BO6),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0fcc00cc0f)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_C5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff0ffff)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_DO6),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_BO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffeefffcfffe)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_CO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.I5(CLBLL_L_X2Y147_SLICE_X1Y147_BO6),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffefffccffee)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y67_I),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_BO6),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_BO6),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_BO6),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000051405140)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_DQ),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_CQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbfffffffa)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_CLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_CO6),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_DO6),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_DO6),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeea4440eeea4440)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aacceef0fafcfe)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000005404)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_CLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeefffe)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BO6),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_BO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7ffffffef)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5454545410101010)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y148_SLICE_X17Y148_D5Q),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0aff0affffff0a)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f2f000002200)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_BLUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_CQ),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I2(CLBLM_L_X16Y152_SLICE_X22Y152_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I5(CLBLM_R_X5Y144_SLICE_X6Y144_A5Q),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffef001000b0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffe)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_CO6),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_BO6),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_AO6),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h005000dc000000cc)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00220022002200f2)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y67_I),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_B5Q),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_L_X12Y148_SLICE_X17Y148_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044000000f400f0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h004400440044f0f4)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_BLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I3(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00f0f0cccc)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffff5fff)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_CO5),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_CO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_DO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc00ccfacc00)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_DLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaffaa00)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_CLUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0a0a0aff080808)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_DO6),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaafc00)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_BO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafffefffe)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_DLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000e000e0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y148_SLICE_X17Y148_DQ),
.I4(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffee00005544)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I4(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_A5Q),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a2a222222222)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_B5Q),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_BO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_CO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I2(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafaeae05050404)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3a3a3a3a3a0a0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbabbba11101110)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcccccccc)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_D5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_AO6),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_D5Q),
.I4(CLBLM_L_X8Y140_SLICE_X11Y140_DO6),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_AO5),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcccccdcc)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_BO6),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_D5Q),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044aaea0040)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_D5Q),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_DO5),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00500050aeae0404)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y148_SLICE_X17Y148_DQ),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0acacacac)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055004400)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_D5Q),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaffaaf0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X15Y144_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_CO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4400000044000000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0a0a0a0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_CLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecf0203cecf0203)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_CO6),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcfefcaa00aa00)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888bb88bb8888)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_BO6),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000f0eef044)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff3c003c)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X15Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080f0000000f)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_BO6),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff504000005040)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc50fffffff0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_DO6),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfebafebafebaeeaa)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_C5Q),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000f000f00)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_A5Q),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfcff505f000)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_C5Q),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_A5Q),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f000afa0afaf)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff040004)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000e000f0000fcfc)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300b8b88888)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_CLUT (
.I0(CLBLM_R_X13Y143_SLICE_X19Y143_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_A5Q),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffccff66)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeecaaa0eeecaaa0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_CO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_DO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8ddddddddddddddd)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_DQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_B5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_B5Q),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002222ff001111)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0faf0eac0eac0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_DQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ddddf0f000ff)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I2(CLBLM_L_X12Y150_SLICE_X16Y150_A5Q),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0609906006099060)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3a0a088008800)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_B5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_B5Q),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f066f066)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_BLUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_DQ),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffb800aa00b8)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_DQ),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_CO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_BO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_DO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0b1a0e4a0e4)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_AO6),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0e4ffffaaff)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00aaaacccc)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_BLUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aaf0aaf0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00000000000000)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_DQ),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff77ffffff)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_CLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020002)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_BLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I2(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_DO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_CO6),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f3fc030c)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_C5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_DO5),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_CO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_DO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50eeee4444)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0faf00a000a00)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0acaca0a0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030ffcc3300)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcceedd33002211)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_DLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_CO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_DO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fc0cf000fc0c)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_C5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefe4454eefe4454)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X13Y142_SLICE_X18Y142_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_BO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_CO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_DO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff005454)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_DLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaefeae54045404)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafcfafc0a0c0a0c)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_BLUT (
.I0(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I4(1'b1),
.I5(CLBLM_L_X12Y147_SLICE_X17Y147_BQ),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbba1110fffa5550)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_DO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddd88888dd8)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_CQ),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I3(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_CO6),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff55f0f0cc44)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_CLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_CQ),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f10101f4f40404)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_CO6),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe54fe54fe54)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_DO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00fa00fa)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_DLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_DQ),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00cc00cc)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_CLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_DQ),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc0f0cf0fc000c)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.I5(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffcc00f000cc)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_BQ),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_CQ),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_CO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffefffffff)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_DO5),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0f5a0e4a0e4)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_CQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_D5Q),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00cfc0cfc0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y143_IOB_X1Y144_I),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfcfcffcccccc)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_BO6),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_CO6),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_DO6),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22fc30fc30)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_DLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_DQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1c0d1c0d1c0d1d1)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_CLUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I5(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3030aaaa3030)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffc0f0c0f0c)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y147_SLICE_X15Y147_D5Q),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_AO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_BO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_CO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8aaa8aa0f000f00)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f50505f0f00000)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_CLUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y147_SLICE_X17Y147_AQ),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5a0a0a0f5a0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfdccec11310020)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I5(CLBLM_L_X8Y148_SLICE_X11Y148_CQ),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_CO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500000000)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_DLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaafe55550054)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff004444ff00f0f0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacffcaaaacffc)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_CO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffaaaa0000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fcfc0c0c)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002222ff003030)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_ALUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_CLUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000010001)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555554500000030)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I4(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_AO5),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a2a0000a2a2888a)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_DLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044555550)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_BO6),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h40f050f0a000a000)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcccccffa0ffa0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.I1(CLBLM_L_X8Y151_SLICE_X11Y151_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_BO6),
.I4(CLBLM_L_X12Y144_SLICE_X17Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_BO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88ffaa5500)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd888888888)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_BO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800880000008000)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f000055565555)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8ffa800a800a8)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_BLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I2(CLBLM_R_X11Y138_SLICE_X15Y138_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f055f011f011)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_ALUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5457a8ab5754aba8)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_CLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_CQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_AO6),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_A5Q),
.I5(CLBLM_R_X11Y138_SLICE_X14Y138_AO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_DO6),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_AO6),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_CO6),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_AO6),
.I5(CLBLM_L_X10Y138_SLICE_X13Y138_CO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc27728dd8)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_AO6),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_A5Q),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_BO6),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I4(CLBLM_R_X13Y142_SLICE_X18Y142_A5Q),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X12Y139_AO6),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22fe02fe02)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_DLUT (
.I0(CLBLM_R_X11Y139_SLICE_X14Y139_DO5),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_C5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4411441100005555)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_DO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000c0ffffff3f)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I2(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_A5Q),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00ba10aa00)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(CLBLM_L_X12Y139_SLICE_X16Y139_BQ),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ff33ff3cffccffc)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_A5Q),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55df55df55105510)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_CLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y138_SLICE_X15Y138_BO6),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a5a533cc)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_BLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_B5Q),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_AO6),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_AO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_AO6),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff84a5b7a5)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_ALUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_AO5),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_AO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00fc00ff)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h050a030305050303)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_AO5),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_CO6),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b888b8b8b888)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_BLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfafa0a0a)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_ALUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_B5Q),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_CO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7fffffff7ffff)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4a0e4a0e4e4e4e4)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfafc0a0c)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_BLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_DO6),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc9cfffff0ff)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_ALUT (
.I0(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I4(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_CO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_CO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110011)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_A5Q),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffcc0000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ec20aaaaa0a0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_CQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I4(CLBLM_L_X12Y142_SLICE_X17Y142_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b888b888b8)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_BO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5f0000ff5c0000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_DO6),
.I3(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h005300a3000300f3)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_A5Q),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.I5(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3f3c0f3)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y143_SLICE_X19Y143_BQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00de12cc00de12)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_ALUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000440044)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_AO6),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y137_SLICE_X12Y137_B5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0a0a0a0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff6c0000006c)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_DO6),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeff1000fe0010)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f4ff000f000f)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c5c00f0a0f0a)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X13Y142_SLICE_X18Y142_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ee22ee22)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_BLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aa0caa0c)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_DLUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_BO5),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_CO6),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaffafaa00040004)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000f000f00)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aa88aa88aa88)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_B5Q),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f044f044)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000a0aff000808)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_CQ),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa003caaaa00cc)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_BLUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_CQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32fe32fe32cc00)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_CQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_BO6),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_CO6),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f111c0c0c000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I5(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f00000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3c0ee22ee22)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaa0aaa0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_CQ),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_AO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h008aaaaa0000aa00)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.I5(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f5f50000ffcc)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_B5Q),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc0037373737)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I3(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee5544faea5040)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.I5(CLBLM_L_X10Y147_SLICE_X13Y147_BO6),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_DO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000faaaa00f0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0a0eeee4444)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f101f404f404)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f50005f5f00500)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a0f0a0f0f0c0c0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_DLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0c5c0cac0ca)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_CLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y147_SLICE_X13Y147_BO6),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0ccccaaaa)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_DQ),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff000f666f000)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_ALUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_DO6),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_BO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_CO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa55aa5a55aa55a)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaf0f03300)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_CLUT (
.I0(CLBLM_R_X13Y142_SLICE_X18Y142_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I3(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafff0aaaaccc0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_BLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff448800004488)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.I3(CLBLM_L_X12Y146_SLICE_X17Y146_CQ),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00020f0d00000f0f)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_CLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_AQ),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf707f808ff0ff000)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_BLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f000f0f07080)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_B5Q),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_CQ),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_CO5),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_AO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_CO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_DO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaaf0f0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000ccacacaca)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fcfc0c0c)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00af05aa00fa50)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_DO6),
.I3(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0d)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_DLUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_AO6),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_CQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.I5(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0000fcdc000a)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c8c8c8c8c8d1c8)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_BLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_ALUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_B5Q),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_BO6),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_CO6),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habeaaabe01400014)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_DO6),
.I5(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f40404fff00f00)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefefa0e0e0e0a)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_DO6),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_AO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbffffffff)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_DLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000200)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_A5Q),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_BLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.I1(CLBLM_L_X12Y148_SLICE_X16Y148_CO6),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0e4a0b1a0e4)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_AO5),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_BO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_CO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_DO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaa5000feaa5400)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaeefa00504450)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404ff0ff000)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I4(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050ccccff00)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_BO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_CO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_DO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaeaffff5040)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeaea40404040)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y146_SLICE_X17Y146_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f00300f3f00300)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y151_SLICE_X18Y151_CQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cfcfc0c0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5454aaaa5454aaa8)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I1(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd8855550505)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I2(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I3(CLBLM_R_X13Y148_SLICE_X19Y148_AQ),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80c0aaff2030aaff)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_BO6),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00d0dddd00d0dddd)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_CO6),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc3333cc33)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h999a9a9999999999)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_CLUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I3(CLBLM_R_X11Y151_SLICE_X14Y151_CO6),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00bf00af00bf00ff)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_BLUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_CO6),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I5(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c5f0c0f4c5f0c0f)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_DO6),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_BQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_BO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9d9d119d1a1bde1b)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fc0cfc0c)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888d8d888888dd8)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_CO6),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h333f333f337f337f)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_DLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_AO5),
.I4(1'b1),
.I5(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05a5a0f3c0ff0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff3100ffff)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AO6),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h333333320000aaaf)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555551ffffffff)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I3(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff040404040)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I3(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X16Y139_AO6),
.Q(CLBLM_L_X12Y139_SLICE_X16Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X16Y139_BO6),
.Q(CLBLM_L_X12Y139_SLICE_X16Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3377337733773377)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_DLUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_DO5),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y141_SLICE_X16Y141_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff1fff00ff1fff00)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_CLUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_DO5),
.I1(CLBLM_L_X12Y141_SLICE_X16Y141_CQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(CLBLM_L_X12Y139_SLICE_X16Y139_BQ),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcccfcccf000f444)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_BLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.I1(CLBLM_R_X13Y150_SLICE_X18Y150_BO6),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_BO6),
.I5(CLBLM_L_X12Y139_SLICE_X16Y139_CO6),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeccfdccfa00f500)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_ALUT (
.I0(CLBLM_L_X12Y139_SLICE_X16Y139_DO6),
.I1(CLBLM_L_X12Y141_SLICE_X16Y141_CQ),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_AQ),
.I3(CLBLM_R_X13Y150_SLICE_X18Y150_BO6),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X17Y139_AO6),
.Q(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X17Y139_BO6),
.Q(CLBLM_L_X12Y139_SLICE_X17Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X17Y139_CO6),
.Q(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X17Y139_DO6),
.Q(CLBLM_L_X12Y139_SLICE_X17Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfafa0000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_DLUT (
.I0(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I2(CLBLM_L_X12Y139_SLICE_X17Y139_DQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0c0f0c0)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_CLUT (
.I0(CLBLM_L_X12Y141_SLICE_X17Y141_CQ),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000cccc)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_BLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaac00c)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_ALUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y148_SLICE_X17Y148_DQ),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X16Y140_AO6),
.Q(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X16Y140_BO6),
.Q(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X16Y140_CO6),
.Q(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a0afa0af)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_DLUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_BO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_DO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefef0f00e0e0000)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_CO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff554400005544)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_BO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddc1110dddc1110)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_AO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_AO6),
.Q(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_BO6),
.Q(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_CO6),
.Q(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011050555440505)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_DLUT (
.I0(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I2(CLBLM_R_X11Y141_SLICE_X14Y141_B5Q),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_DO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0af808f808)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_CO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaabbbb11001111)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_L_X12Y141_SLICE_X17Y141_BQ),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_BO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaa5400feaa5400)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.I2(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I4(CLBLM_L_X12Y142_SLICE_X17Y142_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_AO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X16Y141_BO6),
.Q(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X16Y141_CO5),
.Q(CLBLM_L_X12Y141_SLICE_X16Y141_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X16Y141_AO6),
.Q(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X16Y141_CO6),
.Q(CLBLM_L_X12Y141_SLICE_X16Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_DLUT (
.I0(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.I2(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_DO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afafa0a0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_CLUT (
.I0(CLBLM_L_X12Y139_SLICE_X16Y139_AQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y142_SLICE_X16Y142_A5Q),
.I4(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_CO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc0005050505)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_BO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88d888dd88d8)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I2(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I4(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_AO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X17Y141_AO6),
.Q(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X17Y141_BO6),
.Q(CLBLM_L_X12Y141_SLICE_X17Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X17Y141_CO6),
.Q(CLBLM_L_X12Y141_SLICE_X17Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_DLUT (
.I0(CLBLM_L_X12Y139_SLICE_X17Y139_BQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_AQ),
.I3(CLBLM_L_X12Y141_SLICE_X17Y141_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_DO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a8a8a8a8)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_L_X12Y141_SLICE_X17Y141_CQ),
.I2(CLBLM_L_X12Y139_SLICE_X17Y139_DQ),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_CO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf000f0ccf000)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y141_SLICE_X17Y141_BQ),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_BO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfe0032ccfe0032)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_ALUT (
.I0(CLBLM_L_X12Y141_SLICE_X17Y141_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I4(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_AO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X16Y145_DO6),
.Q(CLBLM_L_X12Y142_SLICE_X16Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X16Y142_AO6),
.Q(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X16Y142_BO6),
.Q(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X16Y142_CO6),
.Q(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff11110000eeee)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_DLUT (
.I0(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DQ),
.I5(CLBLM_R_X13Y142_SLICE_X18Y142_CQ),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_DO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000feaa5400)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X13Y145_SLICE_X18Y145_AQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_CO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0001016868)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_BLUT (
.I0(CLBLM_L_X12Y142_SLICE_X16Y142_DO6),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_DQ),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_B5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_BO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dc10cc00cc00)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.I3(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_AO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X17Y142_AO6),
.Q(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X17Y142_BO6),
.Q(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X17Y142_CO6),
.Q(CLBLM_L_X12Y142_SLICE_X17Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X17Y142_DO6),
.Q(CLBLM_L_X12Y142_SLICE_X17Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeefcfcfccc)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_DLUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_DO6),
.I2(CLBLM_L_X12Y142_SLICE_X17Y142_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_DO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcfc00)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_CLUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_CQ),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_CO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d0c0d0c0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_BO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3e2f3f3f3f3f3)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_ALUT (
.I0(CLBLM_R_X13Y146_SLICE_X18Y146_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_A5Q),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_AO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_BO5),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_CO5),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_AO6),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_BO6),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_CO6),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_A5Q),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_DQ),
.I3(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bbbb8888)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_CLUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X13Y145_SLICE_X18Y145_BQ),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f08888aaaaff00)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_BLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe3332ccdc0010)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_CQ),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X17Y143_AO5),
.Q(CLBLM_L_X12Y143_SLICE_X17Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X17Y143_BO5),
.Q(CLBLM_L_X12Y143_SLICE_X17Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X17Y143_AO6),
.Q(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X17Y143_BO6),
.Q(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X17Y143_CO6),
.Q(CLBLM_L_X12Y143_SLICE_X17Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.Q(CLBLM_L_X12Y143_SLICE_X17Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5e4ffffa0a0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y143_SLICE_X16Y143_B5Q),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_R_X11Y144_SLICE_X15Y144_DO6),
.I5(CLBLM_L_X12Y143_SLICE_X17Y143_DQ),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55550000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y148_SLICE_X17Y148_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaea4040dd88dd88)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I4(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0a0aaee0044)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X13Y142_SLICE_X18Y142_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X17Y144_AO6),
.Q(CLBLM_L_X12Y144_SLICE_X16Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X16Y144_AO6),
.Q(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X16Y144_BO6),
.Q(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X16Y144_DO6),
.Q(CLBLM_L_X12Y144_SLICE_X16Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacac0c0c0c0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4a0cccccc00)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_A5Q),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AQ),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcaff0a00ca000a)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_BLUT (
.I0(CLBLM_R_X13Y145_SLICE_X18Y145_DQ),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fca8fca8)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_AO6),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X16Y144_CO6),
.Q(CLBLM_L_X12Y144_SLICE_X17Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X17Y144_BO6),
.Q(CLBLM_L_X12Y144_SLICE_X17Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X17Y144_CO6),
.Q(CLBLM_L_X12Y144_SLICE_X17Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_DLUT (
.I0(CLBLM_R_X13Y143_SLICE_X19Y143_BQ),
.I1(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.I2(CLBLM_R_X13Y146_SLICE_X19Y146_AQ),
.I3(CLBLM_R_X13Y145_SLICE_X18Y145_DQ),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_DQ),
.I5(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000e0eff000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_CLUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I1(CLBLM_L_X12Y144_SLICE_X17Y144_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X12Y144_SLICE_X17Y144_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20ff33ec20cc00)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_BLUT (
.I0(CLBLM_L_X12Y144_SLICE_X17Y144_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(CLBLM_L_X12Y146_SLICE_X17Y146_BQ),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff0033fffffafa)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_ALUT (
.I0(CLBLM_R_X13Y145_SLICE_X18Y145_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y145_SLICE_X18Y145_CQ),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.Q(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.Q(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X16Y145_CO6),
.Q(CLBLM_L_X12Y145_SLICE_X16Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4a0cccccc00)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_DQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I4(CLBLM_R_X11Y145_SLICE_X15Y145_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005454ff000000)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_CQ),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_AQ),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffccf0c0)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_BLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_B5Q),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd8ddd888d888)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y145_SLICE_X18Y145_DQ),
.I2(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.Q(CLBLM_L_X12Y145_SLICE_X17Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X17Y145_BO6),
.Q(CLBLM_L_X12Y145_SLICE_X17Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.Q(CLBLM_L_X12Y145_SLICE_X17Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X17Y145_DO6),
.Q(CLBLM_L_X12Y145_SLICE_X17Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0cc0000a0cc)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y145_SLICE_X18Y145_BQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafaee50505044)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_CQ),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0f5a0e4e4)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_BQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AQ),
.I3(CLBLM_L_X12Y147_SLICE_X17Y147_BQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeee00000eee0)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_BO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_DO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0fcc00ccf0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_DO5),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e0e01f1f1f1f)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_CLUT (
.I0(CLBLM_R_X13Y145_SLICE_X18Y145_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X13Y145_SLICE_X18Y145_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f4f401010404)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_CO5),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_A5Q),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffee33223322)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_ALUT (
.I0(CLBLM_L_X12Y152_SLICE_X16Y152_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y144_SLICE_X16Y144_A5Q),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_AO6),
.Q(CLBLM_L_X12Y146_SLICE_X17Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_BO6),
.Q(CLBLM_L_X12Y146_SLICE_X17Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.Q(CLBLM_L_X12Y146_SLICE_X17Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4a0cccccc00)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X13Y146_SLICE_X19Y146_AQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000c0c0c0c)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y146_SLICE_X17Y146_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf50d05f8f00800)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_DQ),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33003000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_ALUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y146_SLICE_X17Y146_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_AO6),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_BO6),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_CO6),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f000f000)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00044f0f0ffee)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_CQ),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_AO6),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeee00000eee0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_BLUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_DO6),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeea4440eeea4440)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.I4(CLBLM_R_X13Y148_SLICE_X18Y148_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X17Y147_AO6),
.Q(CLBLM_L_X12Y147_SLICE_X17Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X17Y147_BO6),
.Q(CLBLM_L_X12Y147_SLICE_X17Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X17Y147_CO6),
.Q(CLBLM_L_X12Y147_SLICE_X17Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5550555055554444)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_CQ),
.I2(CLBLM_L_X12Y146_SLICE_X17Y146_AQ),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_DQ),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00a8000000a8)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_CQ),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafc00)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_BLUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_BQ),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccc0aaaaccc0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_DQ),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I2(CLBLM_L_X12Y147_SLICE_X17Y147_AQ),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.Q(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.R(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_CQ),
.Q(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.R(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffafffaf)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_CLUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_BQ),
.I3(CLBLM_R_X13Y147_SLICE_X18Y147_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f000e0e0e0e)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_BLUT (
.I0(CLBLM_L_X12Y149_SLICE_X16Y149_DQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I3(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8bb800f000f0)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_ALUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_DO5),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_AO6),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_BO6),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_CO6),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_DO6),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccf0ccf0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_DLUT (
.I0(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y148_SLICE_X18Y148_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffe0ef000f404)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X12Y148_SLICE_X17Y148_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y150_SLICE_X17Y150_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4e4a0a0a0a0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y147_SLICE_X18Y147_CQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y148_SLICE_X17Y148_BQ),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefff55554555)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X13Y146_SLICE_X18Y146_DO6),
.I5(CLBLM_R_X13Y151_SLICE_X18Y151_CQ),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_AO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_BO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_DO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff00a8a8)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_DO6),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_DQ),
.I3(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa00f0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_CLUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0aaccaaf0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_BLUT (
.I0(CLBLM_L_X12Y146_SLICE_X17Y146_CQ),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaa3330)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_DQ),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I3(CLBLM_L_X12Y150_SLICE_X17Y150_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_AO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_BO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_DO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f20202f2f00200)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I4(CLBLM_L_X12Y148_SLICE_X17Y148_BQ),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_DQ),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff50d8000050d8)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_CLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404ff0ff000)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_BLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_DQ),
.I4(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10dc10ff33cc00)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y150_SLICE_X18Y150_AO5),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y151_SLICE_X19Y151_AO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_BO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_CO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3cff3cff33ff3c)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I2(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I5(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005454ff005151)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_CLUT (
.I0(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfcfc0c0caca)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_CO6),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I5(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f2f2f202020202)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_ALUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_DO6),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X17Y150_AO6),
.Q(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X17Y150_BO6),
.Q(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X17Y150_CO6),
.Q(CLBLM_L_X12Y150_SLICE_X17Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X17Y150_DO6),
.Q(CLBLM_L_X12Y150_SLICE_X17Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1c0d1c0f3f3c0c0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_DLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I3(CLBLM_L_X12Y150_SLICE_X17Y150_DQ),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ee44fa50fa50)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y150_SLICE_X17Y150_CQ),
.I2(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afacafa0a0aca0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I1(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I5(CLBLM_L_X12Y150_SLICE_X17Y150_DQ),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff50ccccff5a)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_ALUT (
.I0(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I2(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y151_SLICE_X17Y151_AO5),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.R(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.R(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.R(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0e0d0f0f0f0f0f)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_DLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I2(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I3(CLBLM_R_X13Y151_SLICE_X18Y151_DO6),
.I4(CLBLM_L_X12Y153_SLICE_X17Y153_CO6),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0d0d0ff0f2f2f0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_CLUT (
.I0(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I2(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3233333333313333)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_BLUT (
.I0(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I2(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I4(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc00dddddddd)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y150_SLICE_X17Y150_DQ),
.Q(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.R(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555fffdffff)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_DLUT (
.I0(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I5(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff001dffff0000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_CLUT (
.I0(CLBLM_R_X13Y151_SLICE_X19Y151_BO6),
.I1(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I2(CLBLM_R_X13Y151_SLICE_X19Y151_CO6),
.I3(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I5(CLBLM_L_X12Y150_SLICE_X17Y150_DQ),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc339c333c)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_BLUT (
.I0(CLBLM_R_X13Y151_SLICE_X19Y151_CO6),
.I1(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.I3(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I4(CLBLM_R_X13Y151_SLICE_X19Y151_BO6),
.I5(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0313ffff00550055)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_ALUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_DO5),
.I2(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I4(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X16Y152_AO6),
.Q(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X16Y152_BO6),
.Q(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000800000a0a0000)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_DLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_CO6),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_DO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaf33333332)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_CLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_CO5),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0efa0afe0efe0e)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_BLUT (
.I0(CLBLM_L_X12Y152_SLICE_X16Y152_DO6),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I5(CLBLM_L_X12Y154_SLICE_X16Y154_BO6),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_BO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfeef00003223)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_ALUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_BO6),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_AO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X17Y152_AO6),
.Q(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X17Y152_BO6),
.Q(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000bbbfffff4440)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_DLUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I1(CLBLM_L_X12Y150_SLICE_X17Y150_CQ),
.I2(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I3(CLBLM_R_X13Y152_SLICE_X18Y152_CO6),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I5(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_DO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5454101054541010)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_CLUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.I2(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I3(1'b1),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_CO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0600000f06)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_CO6),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I2(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y149_SLICE_X13Y149_CQ),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_BO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f0acccc0f0a)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_ALUT (
.I0(CLBLM_L_X12Y152_SLICE_X17Y152_DO6),
.I1(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I2(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_AO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X16Y153_AO6),
.Q(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_DLUT (
.I0(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.I1(CLBLM_L_X12Y153_SLICE_X17Y153_CO6),
.I2(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I4(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I5(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_DO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3000000c70000008)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_CLUT (
.I0(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I5(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_CO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbebeafbebebebebe)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_BLUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I2(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I5(CLBLM_L_X12Y153_SLICE_X16Y153_CO6),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_BO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfc0c0c0cfc0)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_BO6),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_AO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X17Y153_AO6),
.Q(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000100)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_DLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I3(CLBLM_L_X12Y153_SLICE_X17Y153_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_DO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005000400)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_CLUT (
.I0(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I2(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_CO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0780f0ff03c)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_BLUT (
.I0(CLBLM_L_X12Y153_SLICE_X17Y153_DO6),
.I1(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.I2(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.I3(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I5(CLBLM_R_X13Y152_SLICE_X18Y152_DO6),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_BO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfcac0c0cfca)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_ALUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y153_SLICE_X17Y153_BO6),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_AO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X16Y154_AO6),
.Q(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_DO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_CO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h550000038ac3cfc0)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_BLUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I3(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0a0a0afa0a3)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_ALUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I5(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_AO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_DO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_CO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_BO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_AO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X16Y159_DO5),
.O6(CLBLM_L_X12Y159_SLICE_X16Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X16Y159_CO5),
.O6(CLBLM_L_X12Y159_SLICE_X16Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X16Y159_BO5),
.O6(CLBLM_L_X12Y159_SLICE_X16Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_ALUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X16Y159_AO5),
.O6(CLBLM_L_X12Y159_SLICE_X16Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X17Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X17Y159_DO5),
.O6(CLBLM_L_X12Y159_SLICE_X17Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X17Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X17Y159_CO5),
.O6(CLBLM_L_X12Y159_SLICE_X17Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X17Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X17Y159_BO5),
.O6(CLBLM_L_X12Y159_SLICE_X17Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X17Y159_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X17Y159_AO5),
.O6(CLBLM_L_X12Y159_SLICE_X17Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_DO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_CO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_BO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fffffffaa)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(1'b1),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_AO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_DO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_CO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_BO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_AO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_DO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00faf0aa00af0f)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_DO6),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44aa00be14aa00)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_CQ),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_CO6),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff05ff44ff04)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_BLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_DO6),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AO6),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444f5a0f5a0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y127_IOB_X1Y127_I),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_AO5),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffffffff)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000c20002)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_DQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I4(LIOB33_X0Y57_IOB_X0Y58_I),
.I5(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000910080)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(LIOB33_X0Y57_IOB_X0Y57_I),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I5(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000f8f00000)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaffbaffbabababa)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_CLUT (
.I0(CLBLM_R_X3Y144_SLICE_X2Y144_AO6),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdffffeffffff)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111111111111111)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_DLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff2f222f22)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_BLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_DO6),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_DO6),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_CO6),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_DO6),
.I4(CLBLL_L_X4Y145_SLICE_X5Y145_BO6),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_AO6),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdcffffffdcdc)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.I1(CLBLL_L_X2Y146_SLICE_X1Y146_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_BO6),
.I5(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff3dfdfffff)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbffbfffff)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefefeffdfdfdfd)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff101010ff10ff10)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_ALUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I2(LIOB33_X0Y67_IOB_X0Y68_I),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aff0a0aceffcece)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_DLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_B5Q),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeefeffffaafa)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_CLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_AO6),
.I1(CLBLM_L_X16Y152_SLICE_X22Y152_AO6),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_CO6),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000a0000008a88)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_AO6),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffba)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_BO6),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_BO6),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_AO6),
.I5(CLBLL_L_X2Y147_SLICE_X1Y147_AO6),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00eeccfaf0fefc)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_DLUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_DQ),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(CLBLM_L_X16Y152_SLICE_X22Y152_AO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_CLUT (
.I0(CLBLL_L_X2Y147_SLICE_X1Y147_CO6),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_CO6),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_DO6),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_CO6),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BO6),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_ALUT (
.I0(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BO6),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_BO6),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_CO6),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_CO6),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_BO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLM_L_X16Y152_SLICE_X22Y152_AO6),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4f4f4f4fff4f4)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_BLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffffffffff7f)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff0011)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.I1(CLBLL_L_X2Y147_SLICE_X1Y147_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_CO6),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_BO6),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_CO6),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffefffffff)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_AO6),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.I1(CLBLL_L_X2Y147_SLICE_X1Y147_BO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_BO6),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_AO6),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000250fffffeff)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010000000)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.I5(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000f3cc00)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.I2(CLBLL_L_X2Y147_SLICE_X1Y147_BO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffef00200010)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbfffff)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f5f5f1fff5ff)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I2(CLBLM_L_X16Y152_SLICE_X22Y152_AO6),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaeaaaaaa)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_BLUT (
.I0(CLBLM_L_X16Y152_SLICE_X22Y152_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h20200200fffffdff)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffdf00008800)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff0f0f000000)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbfffb)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(1'b1),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_BLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BO5),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_AO5),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffb0000f3f3)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_AO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h050f55ff69966996)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0550cccc0000)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_CO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_BO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff007878)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I3(CLBLM_L_X12Y141_SLICE_X16Y141_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0b1a00000cccc)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_A5Q),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_A5Q),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaaf888f888)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_BLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_A5Q),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555000550050)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_BO5),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_BO6),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_BLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.I1(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc00cc50cc00)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I2(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y139_SLICE_X6Y139_CO6),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_BO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00055ff55ff)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0e0000000e)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_BLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_DO6),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00bb11ba10)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeaaaaa00c00000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_DLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_A5Q),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000001010f000f00)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_CLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_CO6),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0c0f0c0f0c0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5ccffcca0cc00)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_CO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_BO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_DO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfeccde00fa005a)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I3(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0ffc0c0a0a0a0a0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_CO6),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaaaaaf8f88888)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_BLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccf0f000ff)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_ALUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_DO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaafefe54005454)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0eac0faf0eac0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_CLUT (
.I0(CLBLM_L_X12Y143_SLICE_X16Y143_C5Q),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0dff0ff808f000)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4cccc)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_AO5),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_CO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3030aaaa0000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0e4a0e4a0e4a0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cac0c0c0cac0c0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50dddd8888)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_DO5),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_CO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_DO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0aff0ff000)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_B5Q),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4f5e4e4e4e4e4)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f05544)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_BLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ddddd0d0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_BO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_CO5),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_AO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_CO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aaf0fa00aaf0fa)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fa50e4e4e4e4)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_A5Q),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf15fb51f0f00000)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_DQ),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_CQ),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff48c0000048c0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_ALUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_AO6),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff2f3f0f0f)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0fcfc05000c0c)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0fff000c000f0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_DLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_DO6),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_CO6),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_DO6),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_CO6),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_DO6),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_BO6),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3102330033003300)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_CO6),
.I2(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0c0c0c0c0c0c0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacafffff000)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_AO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfddffffcfcc)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_CLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_DO6),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_DO6),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4a0e4f5e4a0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcced00a550505050)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_ALUT (
.I0(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505000037053300)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_DLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff4f4fffffff4)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_CLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_DO6),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fd55ddf0fc00cc)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_BLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.I4(CLBLM_L_X16Y152_SLICE_X22Y152_AO6),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_ALUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_DO6),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_BO6),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_DO6),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_CO6),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h75307530ffff7530)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_DLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_DQ),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44f444f4ffff44f4)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_CLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.I4(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222f2f2ff22fff2)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ccccf0f0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff44fff4)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_DLUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I1(LIOB33_X0Y65_IOB_X0Y66_I),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_DQ),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0caeffff0cae0cae)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_CLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_BQ),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0537003305050000)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_DQ),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888cccca0a0f0f0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffe)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_DLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_AO6),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_CO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_BO6),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000003030ba30)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000a333b000a)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I2(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000a0a33003b0a)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I2(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a0affffff0a)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_DLUT (
.I0(CLBLM_L_X12Y147_SLICE_X17Y147_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.I3(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_BO6),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfe)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_CO6),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_DO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_AO5),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_DO6),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcceefffffcfe)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_BO6),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_AO6),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_AO5),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0c0cccee0cae)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_D5Q),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff5dffffff0c)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_AO6),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_BO6),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000a333b000a)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_CLUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I5(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000d08)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000330050507350)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_DLUT (
.I0(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000b00000008)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h030303ab000000aa)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I4(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_BQ),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffffffffffdff)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000400050000)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3ffffffcffff)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X8Y139_AO6),
.Q(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccf7f7f7f7)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I2(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_AO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ec2000000f0f)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_ALUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I4(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_AO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heece2202ffdf3313)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I5(LIOB33_X0Y53_IOB_X0Y53_I),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcffff)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_D5Q),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_D5Q),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_CLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_D5Q),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_AO6),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffe)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_BO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_BO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff31ffffffff)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I1(LIOB33_X0Y53_IOB_X0Y53_I),
.I2(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_B5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacff0ff000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I4(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffacccc0050)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_BO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_CO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00eeccaa00eecc)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_CQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0c5c0cac0ca)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_B5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff320032ff000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_ALUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1133f1f355fff5ff)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_DLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00005f130000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_CLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I5(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fff88888888)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_BLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000ee88888888)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff5555555555)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5a0e4e4e4e4)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222e2e2e2e2)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003232ff00fafa)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I1(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a000a0000000000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_C5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacc00aaaacc00)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_DQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0caaaaaa00)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y147_SLICE_X15Y147_BQ),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f202f000f000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_ALUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_DO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcac5c0cfcfc0c0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_DLUT (
.I0(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_DQ),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habba0110abba0110)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fef40f000e04)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_DQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafa0000fafa)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_ALUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaafafaaaa)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_DLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_CO6),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I5(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc8888ccc0ccc0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_C5Q),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000ccf0f055cc)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0cac0c5c0ca)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_DO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8dddd8888)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000f000f000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f03300aaaaf0f0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0c0c0c0c0c0c0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_B5Q),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_CQ),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_CO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbb000033330000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_DLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_A5Q),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafaaaa05050000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I5(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f0f005050000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a3aca3ac)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000000000)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_CLUT (
.I0(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_DO6),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc50ffcccc5050)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X9Y145_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y145_SLICE_X9Y145_CO6),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54fe54aa00)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5f5f5e4a0a0a0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3c00aaaacc00)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_BLUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f00ccccf000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbbffbb)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafafa0aca0a0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f0f005050000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ff00f0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_CO5),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_CO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0a0accccff00)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_DLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haeae0404dd88dd88)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0aca0ac)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_DQ),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554555400540054)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_BO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_CO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_DO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff55ccccf050)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_DLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_DQ),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4f5e4a0e4a0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf0f0cccc)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_BLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffe2aa0000e2aa)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_ALUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y151_SLICE_X15Y151_CQ),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_BO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_CO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100000)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_DQ),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00af05fa50)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f44444f4f44444)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_BLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_CO6),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888ddd88888)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I3(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_DO5),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_BO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_CO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_DO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccaaccaa)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_DLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I2(CLBLM_L_X12Y148_SLICE_X17Y148_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00f0f0cccc)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I2(CLBLM_L_X12Y148_SLICE_X17Y148_AQ),
.I3(CLBLM_L_X8Y145_SLICE_X10Y145_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0e4f5e4a0e4)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I2(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc0c80000c0c8)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_ALUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_BO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_CO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_DO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd8ddd888d888)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_A5Q),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_D5Q),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeaefea45404540)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa0c0c)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaaff00)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_BO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_CO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_DO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeaea44444040)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I5(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe0e0ef4f40404)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeaf0c0faeaf0c0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaff00a0a0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_BO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_CO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444044ccccc0cc)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afacafac)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_CLUT (
.I0(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccf00000ccf0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_BQ),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba303055005500)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_CO6),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f00300fcf00c00)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AO6),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_BQ),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hebaa4100faaa5000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AO6),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X14Y138_CO6),
.Q(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44000000f0f0f0b4)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(CLBLM_R_X11Y138_SLICE_X15Y138_DO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I4(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050eaea4040)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_A5Q),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020ffdf000f000f)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_BLUT (
.I0(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f870000ff00)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_ALUT (
.I0(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X15Y138_AO6),
.Q(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff50ff50)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_DLUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_DO6),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000005533a533)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_CLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_A5Q),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_BO5),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I4(CLBLM_R_X11Y138_SLICE_X15Y138_BO5),
.I5(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5556555500ffffff)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I4(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f0bbbb)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y138_SLICE_X15Y138_CO6),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X14Y139_BO6),
.Q(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfdfdffdf0020)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I4(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f0fffff8000ffff)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f011f000f000)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_BLUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_DQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y139_SLICE_X14Y139_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff08f7ffff3333)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I4(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_AO6),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_BO6),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_DQ),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I4(CLBLM_L_X12Y141_SLICE_X17Y141_CQ),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000220fdd0f)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_CLUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_AO5),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_AO5),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_C5Q),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I4(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I5(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf80a08faf80a08)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_BLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f0ccff)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y139_SLICE_X15Y139_CO6),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a00000a05000005)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_DO6),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_A5Q),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0220000001100000)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_CLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_B5Q),
.I1(CLBLM_R_X11Y140_SLICE_X15Y140_CO6),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_AO6),
.I3(CLBLM_L_X12Y141_SLICE_X16Y141_CQ),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_DO6),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0af808f808)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_BLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaa0aaa0a)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_CO6),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_AO6),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ff3cffc3ff3cffc)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.I2(CLBLM_R_X13Y142_SLICE_X18Y142_A5Q),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7d7dffffbebe)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_CQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_DO6),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c53535c5c50535)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_ALUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_CQ),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_BO6),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_DO6),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X14Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X14Y141_BO5),
.Q(CLBLM_R_X11Y141_SLICE_X14Y141_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X14Y141_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X14Y141_BO6),
.Q(CLBLM_R_X11Y141_SLICE_X14Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccc0f0f0cccc)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03030303fc0003ff)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bbbb8888)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffca80000fca8)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_DO6),
.I2(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_BO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005002700af008d)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_CQ),
.I3(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I4(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0123010123012323)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.I2(CLBLM_R_X13Y142_SLICE_X18Y142_A5Q),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.I4(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_A5Q),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05ae04af05ae04)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.I4(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00a8a8)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_DO6),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_AO6),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0050cccc0000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.I3(CLBLM_R_X11Y143_SLICE_X15Y143_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_CLUT (
.I0(CLBLM_L_X12Y144_SLICE_X17Y144_AQ),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00cccc0acc0a)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_BLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_B5Q),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000faaaa00f0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_ALUT (
.I0(CLBLM_R_X13Y145_SLICE_X19Y145_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X15Y142_AO6),
.Q(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X15Y142_CO6),
.Q(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X15Y142_DO6),
.Q(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfebafebafebaeeaa)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_DLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_DQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05af05ab01ab01)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0a0ffcc0000)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_A5Q),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I3(CLBLM_L_X12Y142_SLICE_X17Y142_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ffbb5511)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_CO6),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.Q(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y143_SLICE_X14Y143_BO6),
.Q(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f500d500ff00ff)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_A5Q),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_BQ),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0504040400000000)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(CLBLM_L_X12Y141_SLICE_X16Y141_BO5),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaaaccc0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccccf0a0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffee)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I1(CLBLM_R_X13Y142_SLICE_X18Y142_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DQ),
.I5(CLBLM_L_X12Y143_SLICE_X17Y143_CQ),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffe)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_CLUT (
.I0(CLBLM_L_X12Y143_SLICE_X16Y143_DO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_CQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_A5Q),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_DQ),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_CQ),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.I5(CLBLM_R_X13Y142_SLICE_X18Y142_CQ),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_C5Q),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_DQ),
.I3(CLBLM_R_X11Y143_SLICE_X15Y143_BO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I5(CLBLM_R_X11Y143_SLICE_X15Y143_CO6),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.Q(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.Q(CLBLM_R_X11Y144_SLICE_X14Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000030300000002)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_DLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.I2(CLBLM_L_X12Y141_SLICE_X16Y141_BO5),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafef0f40f000f00)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_CLUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffc0cf505f404)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_BLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00aa00aa)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_CQ),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X15Y144_AO6),
.Q(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.Q(CLBLM_R_X11Y144_SLICE_X15Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbff000003030000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_DLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I1(CLBLM_L_X12Y141_SLICE_X16Y141_A5Q),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefaea55445040)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_DO6),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacaca0cccccc00)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_BLUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y144_SLICE_X15Y144_CQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccff00c0c0)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I2(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X14Y145_BO6),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X14Y145_CO6),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f8f000000000)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacaca0a0acac)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_CLUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88b8888888)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b88b888bb88b888)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_ALUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_AO6),
.Q(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.Q(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_CO6),
.Q(CLBLM_R_X11Y145_SLICE_X15Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_DO6),
.Q(CLBLM_R_X11Y145_SLICE_X15Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffb8b8ffffb888)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fcfcfff0f8f8)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y145_SLICE_X15Y145_CQ),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff060600000606)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_BLUT (
.I0(CLBLM_R_X13Y147_SLICE_X18Y147_CQ),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_BO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_DQ),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0cc0000a0cc)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_BQ),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaaaaaac0000000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1050505000404040)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cacac0c0c0c0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_BLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888b888888b888)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_CO6),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_CO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa00fa00ffcc00cc)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_DLUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_BQ),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_CQ),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habab0101baba1010)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y144_SLICE_X15Y144_BO5),
.I3(1'b1),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I5(CLBLM_R_X11Y148_SLICE_X15Y148_BQ),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f055f0aa)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_BLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y146_SLICE_X17Y146_DO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cfc0cfc0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_CO6),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00df00cc00cca0)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc35aa5cc33aa55)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_CLUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_DO6),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_CQ),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_DO6),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_DQ),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h03030303cfcfcfcf)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555565ffffccff)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_DO5),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_AO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_CO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_DO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10dc10f3f3c0c0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_DQ),
.I3(CLBLM_R_X13Y147_SLICE_X18Y147_CQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01111f0f04444)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffaaf0f0cc88)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_BQ),
.I2(CLBLM_R_X13Y147_SLICE_X18Y147_BQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_CO6),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaccccf0f0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_ALUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_CQ),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_BO6),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000f000f0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aaccaaccaacc)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_DO6),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000c0cff000000)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cac0ff00aa00)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_DQ),
.I1(CLBLM_L_X12Y148_SLICE_X17Y148_D5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y148_SLICE_X16Y148_AO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_BO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_CO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33339393)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_DLUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.I2(CLBLM_R_X11Y150_SLICE_X14Y150_DO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5a0f5a0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_BQ),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0a0a0a0af)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_CO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cacacfc0cfc0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_AO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_AO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_BO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_CO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa5555a955)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_DLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_CO6),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f10401f0f00000)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I4(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f13130f0f0303)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I3(1'b1),
.I4(CLBLM_R_X11Y145_SLICE_X15Y145_CQ),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fe54fa50fe54)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.Q(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.Q(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff1fbf)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_DLUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa5555a595)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_CLUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f0f9f0f00009f0f)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y142_SLICE_X17Y142_CQ),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f004f4f4f004f4f)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X15Y148_DO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f000000000000e0)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_DLUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0a000a000a000a)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_CLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0a00000)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_CO6),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000005050)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X15Y150_AO6),
.Q(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X15Y150_BO6),
.Q(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00f700ff00df)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_CO6),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000010)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_CO6),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffccff000f0c0f)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_CO6),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb7330000b733b733)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_ALUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_DO6),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_AO5),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_BO6),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3ccc39cc33cc33)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_DLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a0f0a005000500)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_CLUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X11Y151_SLICE_X14Y151_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbb8b88bb888b)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_BLUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_CO5),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaeeaafcfcf0f0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_ALUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_DO6),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_DQ),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_BO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_CO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55550000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafa0050aaee0044)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_D5Q),
.I5(CLBLM_L_X12Y152_SLICE_X17Y152_CO6),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4455c4f54455c4f5)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.I1(CLBLM_R_X13Y148_SLICE_X19Y148_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_AO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ffd0fff0f0d0d0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_CO6),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_CO6),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_BO6),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000bb00fc)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_CLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I1(CLBLM_L_X12Y150_SLICE_X17Y150_CQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000aa050f050f)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_BLUT (
.I0(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfa0afa0a)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_ALUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_DO6),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_AO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888888888888)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_DLUT (
.I0(CLBLM_R_X13Y148_SLICE_X19Y148_AQ),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33b0ccff0fbff0f0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_CLUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I1(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_BO5),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_DO6),
.I5(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb300a0007b005a00)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_BLUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I3(CLBLM_L_X12Y152_SLICE_X17Y152_CO6),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_DO5),
.I5(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcffecccc03320000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_ALUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X15Y153_AO6),
.Q(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ff7f0c0c0000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_CLUT (
.I0(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I1(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(CLBLM_L_X12Y152_SLICE_X17Y152_CO5),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010101000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_BLUT (
.I0(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b88b8888b888b)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_DO6),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_CO6),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y140_SLICE_X18Y140_AO6),
.Q(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X18Y140_DO5),
.O6(CLBLM_R_X13Y140_SLICE_X18Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X18Y140_CO5),
.O6(CLBLM_R_X13Y140_SLICE_X18Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X18Y140_BO5),
.O6(CLBLM_R_X13Y140_SLICE_X18Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaaf0ff)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_ALUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_DQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y140_SLICE_X17Y140_DO6),
.O5(CLBLM_R_X13Y140_SLICE_X18Y140_AO5),
.O6(CLBLM_R_X13Y140_SLICE_X18Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_DO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_CO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_BO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y141_SLICE_X18Y141_BO6),
.Q(CLBLM_R_X13Y141_SLICE_X18Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y141_SLICE_X18Y141_AO6),
.Q(CLBLM_R_X13Y141_SLICE_X18Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_DO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000000030000)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(CLBLM_R_X13Y146_SLICE_X18Y146_DO6),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_CO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ea4000003333)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y141_SLICE_X18Y141_A5Q),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I4(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc000c0ffc000c0)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.Q(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_DO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_CO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_BO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaffaaf0aaf0)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_ALUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_AO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y147_SLICE_X18Y147_DO6),
.Q(CLBLM_R_X13Y142_SLICE_X18Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y142_SLICE_X18Y142_AO6),
.Q(CLBLM_R_X13Y142_SLICE_X18Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y142_SLICE_X18Y142_BO6),
.Q(CLBLM_R_X13Y142_SLICE_X18Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y142_SLICE_X18Y142_CO6),
.Q(CLBLM_R_X13Y142_SLICE_X18Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdedeededededdede)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_DLUT (
.I0(CLBLM_R_X13Y146_SLICE_X18Y146_AQ),
.I1(CLBLM_R_X13Y142_SLICE_X18Y142_AQ),
.I2(CLBLM_L_X12Y148_SLICE_X17Y148_CQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y143_SLICE_X18Y143_CO6),
.I5(CLBLM_R_X13Y143_SLICE_X19Y143_CO6),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_DO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055550000)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X13Y142_SLICE_X18Y142_A5Q),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_CO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffb0f0f0f0b)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_BLUT (
.I0(CLBLM_R_X13Y146_SLICE_X18Y146_DO6),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_AQ),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_BO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0aaf0ccf088)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_ALUT (
.I0(CLBLM_R_X13Y142_SLICE_X18Y142_DO6),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_R_X13Y146_SLICE_X18Y146_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_AO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_DO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_CO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_BO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_AO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.Q(CLBLM_R_X13Y143_SLICE_X18Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y143_SLICE_X18Y143_BO6),
.Q(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0ffffffff0ff0)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_CQ),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_CQ),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_AQ),
.I5(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X18Y143_DO5),
.O6(CLBLM_R_X13Y143_SLICE_X18Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cc3c3c3c33c3c)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y143_SLICE_X18Y143_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_CQ),
.I5(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X18Y143_CO5),
.O6(CLBLM_R_X13Y143_SLICE_X18Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haac0aaffaac0aa00)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I1(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(CLBLM_R_X13Y145_SLICE_X19Y145_CQ),
.O5(CLBLM_R_X13Y143_SLICE_X18Y143_BO5),
.O6(CLBLM_R_X13Y143_SLICE_X18Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeff1000fe0010)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X13Y143_SLICE_X18Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X18Y143_AO5),
.O6(CLBLM_R_X13Y143_SLICE_X18Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y143_SLICE_X19Y143_AO6),
.Q(CLBLM_R_X13Y143_SLICE_X19Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y143_SLICE_X19Y143_BO6),
.Q(CLBLM_R_X13Y143_SLICE_X19Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_BQ),
.I2(CLBLM_R_X13Y145_SLICE_X19Y145_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y143_SLICE_X19Y143_AQ),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X19Y143_DO5),
.O6(CLBLM_R_X13Y143_SLICE_X19Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa55aa5a55aa55a)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.O5(CLBLM_R_X13Y143_SLICE_X19Y143_CO5),
.O6(CLBLM_R_X13Y143_SLICE_X19Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaff4055eaaa4000)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y143_SLICE_X19Y143_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I4(CLBLM_R_X13Y146_SLICE_X18Y146_AQ),
.I5(CLBLM_R_X13Y143_SLICE_X19Y143_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X19Y143_BO5),
.O6(CLBLM_R_X13Y143_SLICE_X19Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044aaee0044)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I5(CLBLM_R_X13Y143_SLICE_X19Y143_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X19Y143_AO5),
.O6(CLBLM_R_X13Y143_SLICE_X19Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc30cc33cc33)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y144_SLICE_X17Y144_BQ),
.I2(CLBLM_L_X12Y144_SLICE_X17Y144_AO5),
.I3(CLBLM_L_X12Y146_SLICE_X17Y146_BQ),
.I4(CLBLM_R_X13Y143_SLICE_X19Y143_DO6),
.I5(CLBLM_L_X12Y144_SLICE_X17Y144_DO6),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_DO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddff88aadd558800)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y144_SLICE_X17Y144_BQ),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_CO5),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_BO6),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_CO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fffffeff)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_BLUT (
.I0(CLBLM_R_X13Y143_SLICE_X19Y143_DO6),
.I1(CLBLM_R_X13Y145_SLICE_X18Y145_BQ),
.I2(CLBLM_R_X13Y145_SLICE_X18Y145_CQ),
.I3(CLBLM_L_X12Y144_SLICE_X17Y144_DO6),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_CQ),
.I5(CLBLM_L_X12Y146_SLICE_X17Y146_BQ),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_BO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0201ffffffffffff)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_ALUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_CO5),
.I1(CLBLM_R_X13Y144_SLICE_X19Y144_BO6),
.I2(CLBLM_R_X13Y144_SLICE_X19Y144_AO6),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_DO6),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_AO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff5affaaffa)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_DLUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(CLBLM_R_X13Y146_SLICE_X19Y146_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_DO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_BQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_BQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_CO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffafaffafa)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_BLUT (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_DO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I5(CLBLM_R_X13Y144_SLICE_X19Y144_CO6),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_BO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddffeeffffddffee)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_ALUT (
.I0(CLBLM_R_X13Y145_SLICE_X18Y145_DQ),
.I1(CLBLM_R_X13Y143_SLICE_X18Y143_DO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y145_SLICE_X18Y145_CQ),
.I4(CLBLM_R_X13Y146_SLICE_X18Y146_AQ),
.I5(CLBLM_L_X12Y148_SLICE_X17Y148_CQ),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_AO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y145_SLICE_X18Y145_AO6),
.Q(CLBLM_R_X13Y145_SLICE_X18Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y145_SLICE_X18Y145_BO6),
.Q(CLBLM_R_X13Y145_SLICE_X18Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y145_SLICE_X18Y145_CO6),
.Q(CLBLM_R_X13Y145_SLICE_X18Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y145_SLICE_X18Y145_DO6),
.Q(CLBLM_R_X13Y145_SLICE_X18Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c0c0aaaa)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_DLUT (
.I0(CLBLM_R_X13Y145_SLICE_X19Y145_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y145_SLICE_X18Y145_DQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_DO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d580d580)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I1(CLBLM_R_X13Y145_SLICE_X18Y145_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X13Y146_SLICE_X19Y146_AQ),
.I4(CLBLM_L_X12Y148_SLICE_X17Y148_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_CO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c0c0aaaa)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_BLUT (
.I0(CLBLM_R_X13Y143_SLICE_X19Y143_BQ),
.I1(CLBLM_R_X13Y145_SLICE_X18Y145_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_BO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd8d8ffffd888)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.I2(CLBLM_R_X13Y145_SLICE_X18Y145_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_AO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y145_SLICE_X19Y145_AO6),
.Q(CLBLM_R_X13Y145_SLICE_X19Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y145_SLICE_X19Y145_BO6),
.Q(CLBLM_R_X13Y145_SLICE_X19Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.Q(CLBLM_R_X13Y145_SLICE_X19Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffaaffaa)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_DLUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_DO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ddf055f088f000)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_CQ),
.I2(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_CO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f0fff088f000)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_BQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(CLBLM_R_X13Y145_SLICE_X18Y145_CQ),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_BO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hececccff20200033)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y145_SLICE_X19Y145_AQ),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_AO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y146_SLICE_X18Y146_AO6),
.Q(CLBLM_R_X13Y146_SLICE_X18Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y146_SLICE_X18Y146_CO6),
.Q(CLBLM_R_X13Y146_SLICE_X18Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_DLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_DO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fac8fac8)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_R_X13Y146_SLICE_X18Y146_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_CO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0e2c0ff00aa00)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_BLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X13Y146_SLICE_X18Y146_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_BO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44ee44fa50)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y144_SLICE_X17Y144_CQ),
.I2(CLBLM_R_X13Y146_SLICE_X18Y146_AQ),
.I3(CLBLM_R_X13Y147_SLICE_X18Y147_AQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_AO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.Q(CLBLM_R_X13Y146_SLICE_X19Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_DO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_CO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_BO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8bb888888bb88)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_ALUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y146_SLICE_X19Y146_AQ),
.I3(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_AO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y147_SLICE_X18Y147_AO6),
.Q(CLBLM_R_X13Y147_SLICE_X18Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y147_SLICE_X18Y147_BO6),
.Q(CLBLM_R_X13Y147_SLICE_X18Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y147_SLICE_X18Y147_CO6),
.Q(CLBLM_R_X13Y147_SLICE_X18Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a003030000)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.I2(CLBLM_R_X13Y148_SLICE_X18Y148_BQ),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_A5Q),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_DO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haabb0011bbaa1100)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_R_X13Y146_SLICE_X18Y146_BO5),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_CO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff020c0000020c)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_BLUT (
.I0(CLBLM_R_X13Y148_SLICE_X18Y148_CQ),
.I1(CLBLM_R_X13Y147_SLICE_X18Y147_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I3(CLBLM_R_X13Y147_SLICE_X18Y147_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y144_SLICE_X17Y144_CQ),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_BO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f3f0f3f0)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I2(CLBLM_R_X13Y147_SLICE_X18Y147_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_AO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_DO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_CO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_BO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_DO6),
.Q(CLBLM_R_X13Y148_SLICE_X18Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y148_SLICE_X18Y148_AO6),
.Q(CLBLM_R_X13Y148_SLICE_X18Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y148_SLICE_X18Y148_BO6),
.Q(CLBLM_R_X13Y148_SLICE_X18Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y148_SLICE_X18Y148_CO6),
.Q(CLBLM_R_X13Y148_SLICE_X18Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000a00000002)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I1(CLBLM_R_X13Y148_SLICE_X18Y148_CQ),
.I2(CLBLM_R_X13Y148_SLICE_X18Y148_BQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.I4(CLBLM_R_X13Y147_SLICE_X18Y147_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb51fe54fb51fe54)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y148_SLICE_X18Y148_CQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I4(CLBLM_R_X13Y148_SLICE_X18Y148_DO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_CO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f60006)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_BLUT (
.I0(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.I1(CLBLM_R_X13Y148_SLICE_X18Y148_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.I4(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_BO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffb0f0f0f0b)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_ALUT (
.I0(CLBLM_R_X13Y146_SLICE_X18Y146_DO6),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X13Y148_SLICE_X18Y148_A5Q),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_AO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.Q(CLBLM_R_X13Y148_SLICE_X19Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_DO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_CO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_BO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_AO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.Q(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X18Y149_BO6),
.Q(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_DO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_CO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000044f044f0)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_BLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_BO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0073734040)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_ALUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I2(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I4(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_AO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_DO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_CO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_BO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_AO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_DO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_CO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0f0f0f0f)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_BO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbafa0afa0)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_ALUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y148_SLICE_X18Y148_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_AO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_DO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_CO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_BO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_AO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y151_SLICE_X18Y151_AO6),
.Q(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y151_SLICE_X18Y151_BO6),
.Q(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y151_SLICE_X18Y151_CO6),
.Q(CLBLM_R_X13Y151_SLICE_X18Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040c0c000000000)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_DLUT (
.I0(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I2(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_DO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f8f80c0c0c08)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_CLUT (
.I0(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_CO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0caa0faa0c)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I1(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I2(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_BO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfafbfa51505150)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(1'b1),
.I5(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_AO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_DO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_CLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I1(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I2(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_CO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_BLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I1(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I2(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_BO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccff0fff0f)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_AO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y152_SLICE_X18Y152_AO6),
.Q(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_DLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I3(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y151_SLICE_X18Y151_DO6),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_DO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_CLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I2(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I3(CLBLM_R_X13Y151_SLICE_X18Y151_DO6),
.I4(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I5(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_CO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h85a5c5f5aaaaa0a0)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_BLUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I2(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafabe00005014)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_CO6),
.I2(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I3(CLBLM_R_X13Y152_SLICE_X18Y152_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X13Y148_SLICE_X18Y148_AQ),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_AO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_DO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_CO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_BO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_AO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X15Y144_SLICE_X20Y144_AO6),
.Q(CLBLM_R_X15Y144_SLICE_X20Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X20Y144_DO5),
.O6(CLBLM_R_X15Y144_SLICE_X20Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X20Y144_CO5),
.O6(CLBLM_R_X15Y144_SLICE_X20Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X20Y144_BO5),
.O6(CLBLM_R_X15Y144_SLICE_X20Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0cccc0000)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X15Y144_SLICE_X20Y144_AO5),
.O6(CLBLM_R_X15Y144_SLICE_X20Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X21Y144_DO5),
.O6(CLBLM_R_X15Y144_SLICE_X21Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X21Y144_CO5),
.O6(CLBLM_R_X15Y144_SLICE_X21Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X21Y144_BO5),
.O6(CLBLM_R_X15Y144_SLICE_X21Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X21Y144_AO5),
.O6(CLBLM_R_X15Y144_SLICE_X21Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X15Y151_SLICE_X20Y151_AO6),
.Q(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_DO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_CO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_BO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfffc30303330)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_AO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_DO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_CO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_BO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_AO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y143_SLICE_X56Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y143_SLICE_X56Y143_DO5),
.O6(CLBLM_R_X37Y143_SLICE_X56Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y143_SLICE_X56Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y143_SLICE_X56Y143_CO5),
.O6(CLBLM_R_X37Y143_SLICE_X56Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y143_SLICE_X56Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y143_SLICE_X56Y143_BO5),
.O6(CLBLM_R_X37Y143_SLICE_X56Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300000000)
  ) CLBLM_R_X37Y143_SLICE_X56Y143_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(RIOB33_X105Y119_IOB_X1Y119_I),
.O5(CLBLM_R_X37Y143_SLICE_X56Y143_AO5),
.O6(CLBLM_R_X37Y143_SLICE_X56Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y143_SLICE_X57Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y143_SLICE_X57Y143_DO5),
.O6(CLBLM_R_X37Y143_SLICE_X57Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y143_SLICE_X57Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y143_SLICE_X57Y143_CO5),
.O6(CLBLM_R_X37Y143_SLICE_X57Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y143_SLICE_X57Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y143_SLICE_X57Y143_BO5),
.O6(CLBLM_R_X37Y143_SLICE_X57Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y143_SLICE_X57Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y143_SLICE_X57Y143_AO5),
.O6(CLBLM_R_X37Y143_SLICE_X57Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_DO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_CO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_BO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_AO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_DO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_CO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_BO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00088880000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y139_IOB_X1Y140_I),
.I2(RIOB33_X105Y139_IOB_X1Y139_I),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(RIOB33_X105Y141_IOB_X1Y141_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_AO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffff0f0ffff)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffccccffff)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffff0f0ffff)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I3(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fafafafaf)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(1'b1),
.I4(CLBLM_R_X13Y147_SLICE_X18Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X6Y138_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X0Y135_BO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_AO6),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_BO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_AO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X0Y135_BO5),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X0Y135_AO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_BO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y127_SLICE_X0Y127_AO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y127_SLICE_X0Y127_AO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X12Y143_SLICE_X16Y143_C5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_L_X12Y143_SLICE_X16Y143_CQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X11Y141_SLICE_X14Y141_BQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X10Y137_SLICE_X12Y137_B5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_L_X8Y139_SLICE_X10Y139_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X7Y142_SLICE_X9Y142_B5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X11Y142_SLICE_X14Y142_C5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X4Y140_BQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X4Y140_CQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y141_SLICE_X163Y141_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_R_X103Y141_SLICE_X163Y141_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X12Y159_SLICE_X16Y159_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X0Y135_AO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X37Y143_SLICE_X56Y143_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_R_X13Y145_SLICE_X19Y145_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_L_X12Y147_SLICE_X17Y147_DO6),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X12Y147_SLICE_X17Y147_DO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X12Y148_SLICE_X16Y148_BO6),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X12Y148_SLICE_X16Y148_BO5),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X12Y159_SLICE_X16Y159_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_R_X13Y151_SLICE_X19Y151_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X13Y145_SLICE_X19Y145_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X12Y147_SLICE_X17Y147_DO6),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X12Y147_SLICE_X17Y147_DO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_L_X12Y148_SLICE_X16Y148_BO6),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X12Y148_SLICE_X16Y148_BO5),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_R_X13Y147_SLICE_X18Y147_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_L_X16Y152_SLICE_X22Y152_AO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_L_X16Y152_SLICE_X22Y152_AO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B = CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D = CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_AMUX = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A = CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B = CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C = CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D = CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C = CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D = CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_AMUX = CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_BMUX = CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A = CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B = CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C = CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D = CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A = CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B = CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C = CLBLL_L_X2Y135_SLICE_X0Y135_CO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D = CLBLL_L_X2Y135_SLICE_X0Y135_DO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_AMUX = CLBLL_L_X2Y135_SLICE_X0Y135_AO5;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_BMUX = CLBLL_L_X2Y135_SLICE_X0Y135_BO5;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A = CLBLL_L_X2Y135_SLICE_X1Y135_AO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B = CLBLL_L_X2Y135_SLICE_X1Y135_BO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C = CLBLL_L_X2Y135_SLICE_X1Y135_CO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D = CLBLL_L_X2Y135_SLICE_X1Y135_DO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B = CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C = CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D = CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C = CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D = CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_AMUX = CLBLL_L_X2Y147_SLICE_X0Y147_AO5;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D = CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A = CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B = CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C = CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D = CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_AMUX = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_CMUX = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B = CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C = CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A = CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C = CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_AMUX = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_DMUX = CLBLL_L_X4Y139_SLICE_X4Y139_DO5;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A = CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B = CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C = CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D = CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_AMUX = CLBLL_L_X4Y139_SLICE_X5Y139_AO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_AMUX = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_DMUX = CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B = CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_CMUX = CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_AMUX = CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_AMUX = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CMUX = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CMUX = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A = CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B = CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C = CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D = CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CMUX = CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_BMUX = CLBLL_L_X4Y145_SLICE_X4Y145_B5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CMUX = CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_DMUX = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_AMUX = CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A = CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B = CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_DMUX = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_AMUX = CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A = CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B = CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_AMUX = CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A = CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B = CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A = CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_BMUX = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_AMUX = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A = CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B = CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CMUX = CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A = CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B = CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_AMUX = CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_DMUX = CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A = CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B = CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_BMUX = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B = CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_AMUX = CLBLM_L_X8Y141_SLICE_X10Y141_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_CMUX = CLBLM_L_X8Y141_SLICE_X10Y141_C5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_DMUX = CLBLM_L_X8Y141_SLICE_X10Y141_DO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A = CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_AMUX = CLBLM_L_X8Y141_SLICE_X11Y141_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_AMUX = CLBLM_L_X8Y142_SLICE_X11Y142_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_BMUX = CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_DMUX = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_BMUX = CLBLM_L_X8Y143_SLICE_X10Y143_B5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CMUX = CLBLM_L_X8Y143_SLICE_X10Y143_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_CMUX = CLBLM_L_X8Y143_SLICE_X11Y143_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_DMUX = CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_AMUX = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_CMUX = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A = CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_AMUX = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_CMUX = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A = CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B = CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_DMUX = CLBLM_L_X8Y146_SLICE_X10Y146_D5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A = CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B = CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A = CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A = CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B = CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A = CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B = CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_BMUX = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_DMUX = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A = CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C = CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_DMUX = CLBLM_L_X8Y149_SLICE_X11Y149_DO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_DMUX = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A = CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A = CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D = CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_AMUX = CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_BMUX = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A = CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_AMUX = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_DMUX = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_BMUX = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_CMUX = CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_DMUX = CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A = CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A = CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A = CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C = CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_CMUX = CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A = CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B = CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_AMUX = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_BMUX = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A = CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B = CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_AMUX = CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_AMUX = CLBLM_L_X10Y141_SLICE_X12Y141_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_BMUX = CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A = CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_AMUX = CLBLM_L_X10Y142_SLICE_X13Y142_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_BMUX = CLBLM_L_X10Y142_SLICE_X13Y142_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CMUX = CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_DMUX = CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_AMUX = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CMUX = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_BMUX = CLBLM_L_X10Y144_SLICE_X12Y144_B5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_DMUX = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_BMUX = CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_CMUX = CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CMUX = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_BMUX = CLBLM_L_X10Y145_SLICE_X13Y145_B5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_DMUX = CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B = CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C = CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CMUX = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A = CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CMUX = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A = CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A = CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B = CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A = CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A = CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CMUX = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A = CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C = CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_CMUX = CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_AMUX = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A = CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B = CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C = CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A = CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_AMUX = CLBLM_L_X10Y152_SLICE_X13Y152_AO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B = CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C = CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D = CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C = CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A = CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B = CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C = CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D = CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_DMUX = CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A = CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B = CLBLM_L_X12Y140_SLICE_X17Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A = CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B = CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C = CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D = CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_AMUX = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_BMUX = CLBLM_L_X12Y141_SLICE_X16Y141_BO5;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_CMUX = CLBLM_L_X12Y141_SLICE_X16Y141_C5Q;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A = CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B = CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C = CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A = CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B = CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C = CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D = CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_AMUX = CLBLM_L_X12Y142_SLICE_X16Y142_A5Q;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A = CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B = CLBLM_L_X12Y142_SLICE_X17Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C = CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B = CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C = CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_BMUX = CLBLM_L_X12Y143_SLICE_X16Y143_B5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_CMUX = CLBLM_L_X12Y143_SLICE_X16Y143_C5Q;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A = CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B = CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C = CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_AMUX = CLBLM_L_X12Y143_SLICE_X17Y143_A5Q;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_BMUX = CLBLM_L_X12Y143_SLICE_X17Y143_B5Q;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B = CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_AMUX = CLBLM_L_X12Y144_SLICE_X16Y144_A5Q;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_CMUX = CLBLM_L_X12Y144_SLICE_X16Y144_CO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A = CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B = CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C = CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D = CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_AMUX = CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_DMUX = CLBLM_L_X12Y145_SLICE_X16Y145_DO5;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_AMUX = CLBLM_L_X12Y146_SLICE_X16Y146_A5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_CMUX = CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A = CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B = CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_DMUX = CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A = CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B = CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C = CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B = CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C = CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_DMUX = CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D = CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_AMUX = CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_BMUX = CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B = CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C = CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D = CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_DMUX = CLBLM_L_X12Y148_SLICE_X17Y148_D5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A = CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A = CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B = CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C = CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_AMUX = CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_BMUX = CLBLM_L_X12Y150_SLICE_X16Y150_B5Q;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A = CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B = CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C = CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D = CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A = CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_AMUX = CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_DMUX = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B = CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_AMUX = CLBLM_L_X12Y151_SLICE_X17Y151_AO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A = CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B = CLBLM_L_X12Y152_SLICE_X16Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_CMUX = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_DMUX = CLBLM_L_X12Y152_SLICE_X16Y152_DO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A = CLBLM_L_X12Y152_SLICE_X17Y152_AO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B = CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D = CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_CMUX = CLBLM_L_X12Y152_SLICE_X17Y152_CO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A = CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B = CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C = CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A = CLBLM_L_X12Y153_SLICE_X17Y153_AO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B = CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A = CLBLM_L_X12Y154_SLICE_X16Y154_AO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B = CLBLM_L_X12Y154_SLICE_X16Y154_BO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C = CLBLM_L_X12Y154_SLICE_X16Y154_CO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D = CLBLM_L_X12Y154_SLICE_X16Y154_DO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_BMUX = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A = CLBLM_L_X12Y154_SLICE_X17Y154_AO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B = CLBLM_L_X12Y154_SLICE_X17Y154_BO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C = CLBLM_L_X12Y154_SLICE_X17Y154_CO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D = CLBLM_L_X12Y154_SLICE_X17Y154_DO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B = CLBLM_L_X12Y159_SLICE_X16Y159_BO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C = CLBLM_L_X12Y159_SLICE_X16Y159_CO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D = CLBLM_L_X12Y159_SLICE_X16Y159_DO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A = CLBLM_L_X12Y159_SLICE_X17Y159_AO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B = CLBLM_L_X12Y159_SLICE_X17Y159_BO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C = CLBLM_L_X12Y159_SLICE_X17Y159_CO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D = CLBLM_L_X12Y159_SLICE_X17Y159_DO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B = CLBLM_L_X16Y152_SLICE_X22Y152_BO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C = CLBLM_L_X16Y152_SLICE_X22Y152_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D = CLBLM_L_X16Y152_SLICE_X22Y152_DO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_AMUX = CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A = CLBLM_L_X16Y152_SLICE_X23Y152_AO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B = CLBLM_L_X16Y152_SLICE_X23Y152_BO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C = CLBLM_L_X16Y152_SLICE_X23Y152_CO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D = CLBLM_L_X16Y152_SLICE_X23Y152_DO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_AMUX = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A = CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A = CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C = CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_AMUX = CLBLM_R_X3Y144_SLICE_X3Y144_AO5;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B = CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C = CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_AMUX = CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A = CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_AMUX = CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_BMUX = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_CMUX = CLBLM_R_X3Y146_SLICE_X2Y146_CO5;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A = CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B = CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C = CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D = CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_AMUX = CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C = CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B = CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_AMUX = CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A = CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_AMUX = CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_AMUX = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_AMUX = CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_CMUX = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_AMUX = CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_BMUX = CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C = CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_AMUX = CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A = CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A = CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_BMUX = CLBLM_R_X5Y139_SLICE_X6Y139_BO5;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A = CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B = CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A = CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B = CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_AMUX = CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CMUX = CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_BMUX = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CMUX = CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_DMUX = CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CMUX = CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_AMUX = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_BMUX = CLBLM_R_X5Y143_SLICE_X6Y143_B5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CMUX = CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A = CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_AMUX = CLBLM_R_X5Y144_SLICE_X6Y144_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A = CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C = CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_DMUX = CLBLM_R_X5Y144_SLICE_X7Y144_D5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A = CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B = CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C = CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_AMUX = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_BMUX = CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_CMUX = CLBLM_R_X5Y145_SLICE_X6Y145_C5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A = CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B = CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_AMUX = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CMUX = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A = CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B = CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_AMUX = CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B = CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A = CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_AMUX = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_DMUX = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A = CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B = CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A = CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B = CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C = CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_AMUX = CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B = CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D = CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_AMUX = CLBLM_R_X5Y150_SLICE_X6Y150_AO5;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A = CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B = CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C = CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D = CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_AMUX = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A = CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_AMUX = CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_AMUX = CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A = CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B = CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C = CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_AMUX = CLBLM_R_X7Y140_SLICE_X9Y140_AO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A = CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AMUX = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_BMUX = CLBLM_R_X7Y141_SLICE_X8Y141_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_AMUX = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_BMUX = CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_BMUX = CLBLM_R_X7Y142_SLICE_X9Y142_B5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A = CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_AMUX = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_BMUX = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A = CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CMUX = CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_BMUX = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C = CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_DMUX = CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A = CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A = CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CMUX = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A = CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B = CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A = CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B = CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C = CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_DMUX = CLBLM_R_X7Y148_SLICE_X9Y148_D5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A = CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B = CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A = CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A = CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B = CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_AMUX = CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_DMUX = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B = CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A = CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B = CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C = CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B = CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_AMUX = CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_BMUX = CLBLM_R_X11Y138_SLICE_X14Y138_BO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_DMUX = CLBLM_R_X11Y138_SLICE_X14Y138_DO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A = CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_BMUX = CLBLM_R_X11Y138_SLICE_X15Y138_BO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B = CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_AMUX = CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CMUX = CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_DMUX = CLBLM_R_X11Y139_SLICE_X14Y139_DO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A = CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B = CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D = CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A = CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B = CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_AMUX = CLBLM_R_X11Y141_SLICE_X14Y141_A5Q;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_BMUX = CLBLM_R_X11Y141_SLICE_X14Y141_B5Q;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CMUX = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_DMUX = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A = CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B = CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C = CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_BMUX = CLBLM_R_X11Y142_SLICE_X14Y142_B5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CMUX = CLBLM_R_X11Y142_SLICE_X14Y142_C5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A = CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B = CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C = CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D = CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_BMUX = CLBLM_R_X11Y142_SLICE_X15Y142_BO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_CMUX = CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_BMUX = CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A = CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D = CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_CMUX = CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_DMUX = CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_DMUX = CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_AMUX = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_BMUX = CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_CMUX = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_DMUX = CLBLM_R_X11Y147_SLICE_X15Y147_D5Q;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_AMUX = CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_AMUX = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_AMUX = CLBLM_R_X11Y149_SLICE_X14Y149_A5Q;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_AMUX = CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_BMUX = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_CMUX = CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B = CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_AMUX = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CMUX = CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A = CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B = CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D = CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B = CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C = CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_BMUX = CLBLM_R_X11Y152_SLICE_X14Y152_BO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A = CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C = CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D = CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A = CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_BMUX = CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_CMUX = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A = CLBLM_R_X13Y140_SLICE_X18Y140_AO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B = CLBLM_R_X13Y140_SLICE_X18Y140_BO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C = CLBLM_R_X13Y140_SLICE_X18Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D = CLBLM_R_X13Y140_SLICE_X18Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A = CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B = CLBLM_R_X13Y140_SLICE_X19Y140_BO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C = CLBLM_R_X13Y140_SLICE_X19Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D = CLBLM_R_X13Y140_SLICE_X19Y140_DO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A = CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D = CLBLM_R_X13Y141_SLICE_X18Y141_DO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_AMUX = CLBLM_R_X13Y141_SLICE_X18Y141_A5Q;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_BMUX = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A = CLBLM_R_X13Y141_SLICE_X19Y141_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B = CLBLM_R_X13Y141_SLICE_X19Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C = CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D = CLBLM_R_X13Y141_SLICE_X19Y141_DO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B = CLBLM_R_X13Y142_SLICE_X18Y142_BO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C = CLBLM_R_X13Y142_SLICE_X18Y142_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D = CLBLM_R_X13Y142_SLICE_X18Y142_DO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_AMUX = CLBLM_R_X13Y142_SLICE_X18Y142_A5Q;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A = CLBLM_R_X13Y142_SLICE_X19Y142_AO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B = CLBLM_R_X13Y142_SLICE_X19Y142_BO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C = CLBLM_R_X13Y142_SLICE_X19Y142_CO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D = CLBLM_R_X13Y142_SLICE_X19Y142_DO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B = CLBLM_R_X13Y143_SLICE_X18Y143_BO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C = CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D = CLBLM_R_X13Y143_SLICE_X18Y143_DO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A = CLBLM_R_X13Y143_SLICE_X19Y143_AO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B = CLBLM_R_X13Y143_SLICE_X19Y143_BO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C = CLBLM_R_X13Y143_SLICE_X19Y143_CO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D = CLBLM_R_X13Y143_SLICE_X19Y143_DO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_CMUX = CLBLM_R_X13Y143_SLICE_X19Y143_CO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B = CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D = CLBLM_R_X13Y144_SLICE_X18Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_DMUX = CLBLM_R_X13Y144_SLICE_X18Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A = CLBLM_R_X13Y144_SLICE_X19Y144_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B = CLBLM_R_X13Y144_SLICE_X19Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C = CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D = CLBLM_R_X13Y144_SLICE_X19Y144_DO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A = CLBLM_R_X13Y145_SLICE_X18Y145_AO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B = CLBLM_R_X13Y145_SLICE_X18Y145_BO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C = CLBLM_R_X13Y145_SLICE_X18Y145_CO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D = CLBLM_R_X13Y145_SLICE_X18Y145_DO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A = CLBLM_R_X13Y145_SLICE_X19Y145_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B = CLBLM_R_X13Y145_SLICE_X19Y145_BO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A = CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C = CLBLM_R_X13Y146_SLICE_X18Y146_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D = CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_BMUX = CLBLM_R_X13Y146_SLICE_X18Y146_BO5;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B = CLBLM_R_X13Y146_SLICE_X19Y146_BO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C = CLBLM_R_X13Y146_SLICE_X19Y146_CO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D = CLBLM_R_X13Y146_SLICE_X19Y146_DO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A = CLBLM_R_X13Y147_SLICE_X18Y147_AO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B = CLBLM_R_X13Y147_SLICE_X18Y147_BO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C = CLBLM_R_X13Y147_SLICE_X18Y147_CO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D = CLBLM_R_X13Y147_SLICE_X18Y147_DO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_DMUX = CLBLM_R_X13Y147_SLICE_X18Y147_DO5;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A = CLBLM_R_X13Y147_SLICE_X19Y147_AO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C = CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D = CLBLM_R_X13Y147_SLICE_X19Y147_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A = CLBLM_R_X13Y148_SLICE_X18Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B = CLBLM_R_X13Y148_SLICE_X18Y148_BO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C = CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D = CLBLM_R_X13Y148_SLICE_X18Y148_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_AMUX = CLBLM_R_X13Y148_SLICE_X18Y148_A5Q;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_DMUX = CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A = CLBLM_R_X13Y148_SLICE_X19Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B = CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C = CLBLM_R_X13Y148_SLICE_X19Y148_CO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D = CLBLM_R_X13Y148_SLICE_X19Y148_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B = CLBLM_R_X13Y149_SLICE_X18Y149_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C = CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D = CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A = CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B = CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C = CLBLM_R_X13Y149_SLICE_X19Y149_CO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D = CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C = CLBLM_R_X13Y150_SLICE_X18Y150_CO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D = CLBLM_R_X13Y150_SLICE_X18Y150_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_AMUX = CLBLM_R_X13Y150_SLICE_X18Y150_AO5;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A = CLBLM_R_X13Y150_SLICE_X19Y150_AO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B = CLBLM_R_X13Y150_SLICE_X19Y150_BO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C = CLBLM_R_X13Y150_SLICE_X19Y150_CO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D = CLBLM_R_X13Y150_SLICE_X19Y150_DO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A = CLBLM_R_X13Y151_SLICE_X18Y151_AO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B = CLBLM_R_X13Y151_SLICE_X18Y151_BO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C = CLBLM_R_X13Y151_SLICE_X18Y151_CO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D = CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A = CLBLM_R_X13Y151_SLICE_X19Y151_AO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B = CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C = CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D = CLBLM_R_X13Y151_SLICE_X19Y151_DO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_AMUX = CLBLM_R_X13Y151_SLICE_X19Y151_AO5;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A = CLBLM_R_X13Y152_SLICE_X18Y152_AO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B = CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C = CLBLM_R_X13Y152_SLICE_X18Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D = CLBLM_R_X13Y152_SLICE_X18Y152_DO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_BMUX = CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A = CLBLM_R_X13Y152_SLICE_X19Y152_AO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B = CLBLM_R_X13Y152_SLICE_X19Y152_BO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C = CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D = CLBLM_R_X13Y152_SLICE_X19Y152_DO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A = CLBLM_R_X15Y144_SLICE_X20Y144_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B = CLBLM_R_X15Y144_SLICE_X20Y144_BO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D = CLBLM_R_X15Y144_SLICE_X20Y144_DO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D = CLBLM_R_X15Y144_SLICE_X21Y144_DO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A = CLBLM_R_X15Y151_SLICE_X20Y151_AO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B = CLBLM_R_X15Y151_SLICE_X20Y151_BO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C = CLBLM_R_X15Y151_SLICE_X20Y151_CO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A = CLBLM_R_X15Y151_SLICE_X21Y151_AO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B = CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C = CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_A = CLBLM_R_X37Y143_SLICE_X56Y143_AO6;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_B = CLBLM_R_X37Y143_SLICE_X56Y143_BO6;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_C = CLBLM_R_X37Y143_SLICE_X56Y143_CO6;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_D = CLBLM_R_X37Y143_SLICE_X56Y143_DO6;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_A = CLBLM_R_X37Y143_SLICE_X57Y143_AO6;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_B = CLBLM_R_X37Y143_SLICE_X57Y143_BO6;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_C = CLBLM_R_X37Y143_SLICE_X57Y143_CO6;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_D = CLBLM_R_X37Y143_SLICE_X57Y143_DO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A = CLBLM_R_X103Y141_SLICE_X162Y141_AO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B = CLBLM_R_X103Y141_SLICE_X162Y141_BO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C = CLBLM_R_X103Y141_SLICE_X162Y141_CO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D = CLBLM_R_X103Y141_SLICE_X162Y141_DO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B = CLBLM_R_X103Y141_SLICE_X163Y141_BO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C = CLBLM_R_X103Y141_SLICE_X163Y141_CO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D = CLBLM_R_X103Y141_SLICE_X163Y141_DO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_AMUX = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_AMUX = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A = CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B = CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C = CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D = CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B = CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C = CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D = CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_AMUX = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y135_SLICE_X0Y135_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y135_SLICE_X0Y135_BO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X12Y143_SLICE_X16Y143_C5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X7Y142_SLICE_X9Y142_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X4Y140_SLICE_X4Y140_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X11Y142_SLICE_X14Y142_C5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_R_X13Y151_SLICE_X19Y151_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_R_X13Y147_SLICE_X18Y147_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X37Y143_SLICE_X56Y143_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B1 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B2 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B3 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B4 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C2 = CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C3 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C5 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C6 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D3 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D5 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D6 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A1 = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A2 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A3 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A4 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B2 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B3 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B4 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B6 = CLBLM_L_X12Y142_SLICE_X17Y142_CQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A3 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A4 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A5 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C1 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C2 = CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C3 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D1 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D3 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D4 = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A5 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B3 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B4 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B5 = CLBLM_R_X11Y145_SLICE_X15Y145_CQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B6 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_AX = CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A3 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D2 = CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D3 = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D4 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D5 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D6 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C2 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D4 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A2 = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A5 = CLBLM_R_X13Y142_SLICE_X18Y142_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B2 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B4 = CLBLM_L_X8Y141_SLICE_X10Y141_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C3 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C1 = CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C2 = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C4 = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C5 = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C6 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D1 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D4 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D5 = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A3 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A4 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B1 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B2 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B6 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C4 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C6 = CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D2 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D3 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D4 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D5 = CLBLM_L_X12Y150_SLICE_X16Y150_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A1 = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A2 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A3 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A4 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A5 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B1 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B2 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B4 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B5 = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B6 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A1 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A3 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A4 = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A5 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C1 = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C2 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C3 = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B2 = CLBLM_R_X5Y144_SLICE_X7Y144_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B3 = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B5 = CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B6 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D1 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C1 = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C2 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C3 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C4 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C5 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C6 = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D3 = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D4 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A1 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A2 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A3 = CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A4 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A5 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D4 = CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D6 = CLBLM_R_X7Y148_SLICE_X9Y148_D5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B2 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B3 = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B4 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B5 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A4 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A5 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C1 = CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A6 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C1 = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C2 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C3 = CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D1 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D2 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D4 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D5 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D6 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D4 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A2 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A3 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A4 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A5 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A6 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_SR = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B2 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B4 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B5 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B6 = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C1 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C2 = CLBLM_L_X8Y147_SLICE_X11Y147_CQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C3 = CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C4 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C6 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D2 = CLBLM_L_X8Y147_SLICE_X11Y147_CQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D3 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D4 = CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D6 = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A2 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A3 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A4 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A5 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A6 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B1 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B2 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B4 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B6 = CLBLM_L_X12Y147_SLICE_X17Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C2 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C6 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D1 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D2 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D3 = CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D4 = CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D6 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_BX = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A1 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A2 = CLBLM_R_X13Y148_SLICE_X19Y148_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A3 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A5 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C1 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B3 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B5 = CLBLM_R_X7Y148_SLICE_X9Y148_D5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B6 = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C3 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A1 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A3 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C2 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B1 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B2 = CLBLM_R_X7Y141_SLICE_X8Y141_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B6 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C2 = CLBLM_R_X7Y141_SLICE_X9Y141_CQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C4 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C5 = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A1 = CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A3 = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A4 = CLBLM_L_X10Y149_SLICE_X13Y149_DQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B1 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B3 = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B4 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A2 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C4 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AX = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B1 = CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B2 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B5 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D1 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D2 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C1 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C2 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C3 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C5 = CLBLM_R_X7Y141_SLICE_X8Y141_B5Q;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D2 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D3 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D4 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D3 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D4 = CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A2 = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A3 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A4 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B2 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B4 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B5 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C2 = CLBLM_L_X8Y148_SLICE_X11Y148_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C3 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C4 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C6 = CLBLM_R_X5Y144_SLICE_X7Y144_D5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D3 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D4 = CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D5 = CLBLM_L_X8Y149_SLICE_X11Y149_DO5;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D6 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A2 = CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A3 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A6 = CLBLM_L_X8Y149_SLICE_X10Y149_CQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B4 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B5 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B6 = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C1 = CLBLM_L_X8Y149_SLICE_X10Y149_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C2 = CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C4 = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C5 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D1 = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D2 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D3 = CLBLM_L_X8Y148_SLICE_X10Y148_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D4 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C6 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A1 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A3 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A4 = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B1 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B2 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B3 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B4 = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B5 = CLBLM_L_X12Y152_SLICE_X16Y152_DO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B6 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D2 = CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A1 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A2 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_C5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A6 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C1 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C2 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C3 = CLBLM_R_X11Y152_SLICE_X14Y152_BO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B5 = CLBLM_L_X8Y145_SLICE_X10Y145_DQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D5 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D6 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C2 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C6 = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A1 = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A2 = CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A4 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D4 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D6 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A6 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B1 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A4 = CLBLM_L_X10Y143_SLICE_X13Y143_CQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A3 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A4 = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C1 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C2 = CLBLM_L_X12Y150_SLICE_X17Y150_CQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B1 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B3 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B4 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D1 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D2 = CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C1 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C3 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C4 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C5 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C6 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D3 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D4 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D6 = CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B1 = CLBLM_L_X12Y147_SLICE_X16Y147_CQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D1 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D2 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B2 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D3 = CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D4 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D5 = CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D6 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B3 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B4 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B6 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C5 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C4 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A3 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A4 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A5 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A6 = CLBLM_L_X8Y148_SLICE_X11Y148_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B5 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C4 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C1 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C5 = CLBLM_L_X12Y147_SLICE_X17Y147_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C6 = CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C5 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D4 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D2 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A2 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A4 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A6 = CLBLM_R_X11Y147_SLICE_X15Y147_D5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B2 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B3 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C1 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C3 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C4 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C5 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C6 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D3 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D1 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D3 = CLBLM_L_X8Y149_SLICE_X10Y149_DQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D4 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D4 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A1 = CLBLM_R_X7Y147_SLICE_X9Y147_DQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A5 = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A6 = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B1 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B4 = CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B5 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A1 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C1 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C2 = CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B4 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B6 = CLBLM_R_X7Y143_SLICE_X9Y143_DQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C3 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C4 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C5 = CLBLM_R_X7Y142_SLICE_X9Y142_B5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D1 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D2 = CLBLM_R_X13Y145_SLICE_X19Y145_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D4 = CLBLM_R_X7Y143_SLICE_X9Y143_DQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D6 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A1 = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A4 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A5 = CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A6 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_AX = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B2 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B4 = CLBLM_R_X11Y147_SLICE_X15Y147_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B5 = CLBLM_L_X10Y142_SLICE_X13Y142_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C1 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C2 = CLBLM_L_X10Y143_SLICE_X13Y143_DQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_C5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D3 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D4 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D6 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A1 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A4 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A6 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B2 = CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C1 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C6 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A2 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A4 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B1 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B3 = CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B4 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B6 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C2 = CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C3 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C4 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C5 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C6 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D1 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D5 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D6 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A1 = CLBLM_R_X5Y143_SLICE_X6Y143_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A2 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A4 = CLBLM_R_X7Y141_SLICE_X9Y141_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A5 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A6 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B1 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B4 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C3 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C6 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D2 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D3 = CLBLM_R_X7Y144_SLICE_X9Y144_DQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D6 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A1 = CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A5 = CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B2 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B3 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C1 = CLBLM_L_X8Y143_SLICE_X11Y143_C5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C3 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C4 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D1 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D4 = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D5 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D6 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A2 = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A4 = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A5 = CLBLM_L_X12Y144_SLICE_X17Y144_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D4 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D5 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B1 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B2 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B3 = CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B4 = CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B5 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B6 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C3 = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C4 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C5 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D1 = CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D2 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D4 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D5 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D6 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A3 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A4 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A5 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B1 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B2 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B4 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B5 = CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C1 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C3 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C4 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C5 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C6 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D4 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A2 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A3 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A4 = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A6 = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B2 = CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B3 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B4 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B5 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B6 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C1 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C2 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C3 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C4 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C5 = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C6 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D1 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D2 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D3 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A1 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A4 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B5 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B6 = CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C5 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C6 = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D1 = CLBLM_L_X12Y144_SLICE_X16Y144_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D2 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D4 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B2 = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C4 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B1 = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D4 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C1 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A1 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A3 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A4 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A5 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C3 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B5 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B6 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C1 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C2 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C4 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C5 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C6 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D1 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D2 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D4 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A2 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A4 = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A6 = CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B1 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B2 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B4 = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B6 = CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C2 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C3 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C4 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C5 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C6 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D2 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D3 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D4 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D4 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D4 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A6 = CLBLM_R_X13Y148_SLICE_X18Y148_A5Q;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C5 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B4 = CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B5 = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B6 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A1 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A2 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A6 = CLBLM_R_X11Y151_SLICE_X15Y151_CQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D2 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B1 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B2 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B3 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B4 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B6 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C2 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C3 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C4 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C5 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C6 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D5 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C4 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D6 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C5 = CLBLM_R_X13Y148_SLICE_X18Y148_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D1 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D2 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D3 = CLBLM_R_X7Y147_SLICE_X9Y147_DQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D4 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D6 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A1 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A3 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A6 = CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A5 = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B4 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B5 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B6 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C2 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C4 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D1 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D2 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D4 = CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D6 = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D1 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D2 = CLBLM_R_X13Y148_SLICE_X18Y148_CQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D3 = CLBLM_R_X13Y148_SLICE_X18Y148_BQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D4 = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B3 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A2 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A3 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A4 = CLBLM_R_X3Y146_SLICE_X2Y146_CO5;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B2 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B3 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B4 = CLBLM_R_X3Y146_SLICE_X2Y146_CO5;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B5 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C2 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C3 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C4 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C5 = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C6 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A2 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A3 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A5 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A1 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A3 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A6 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B2 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B3 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B4 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B5 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A4 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C3 = CLBLM_L_X12Y148_SLICE_X17Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C4 = CLBLM_L_X8Y145_SLICE_X10Y145_DQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B4 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D1 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A1 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A5 = CLBLM_L_X12Y150_SLICE_X16Y150_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B1 = CLBLM_R_X5Y139_SLICE_X6Y139_BO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B2 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B3 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B4 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B5 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B6 = CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C4 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A1 = CLBLL_L_X2Y147_SLICE_X0Y147_AO5;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A2 = CLBLM_R_X5Y143_SLICE_X6Y143_B5Q;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A3 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A6 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B3 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C4 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y135_SLICE_X0Y135_AO5;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y135_SLICE_X0Y135_BO5;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A2 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A4 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A6 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B2 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B4 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B5 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A1 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A3 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A4 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A5 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C1 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C2 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B1 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B3 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B4 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C4 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D1 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D3 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D4 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D5 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A1 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A2 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A4 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B1 = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B2 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B5 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C1 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C2 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C3 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C4 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C5 = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D6 = CLBLM_R_X7Y148_SLICE_X9Y148_D5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D4 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C3 = CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C4 = CLBLM_L_X12Y141_SLICE_X16Y141_CQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D4 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D5 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D1 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B2 = CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B3 = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B4 = CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D6 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A2 = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A3 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A5 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B2 = CLBLM_R_X7Y150_SLICE_X9Y150_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B3 = CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B4 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B6 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C1 = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C2 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C4 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D4 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D5 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A2 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A4 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B2 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B4 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C2 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C4 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D2 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D4 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D2 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D2 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D3 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D4 = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D5 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D3 = CLBLM_L_X12Y148_SLICE_X17Y148_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D6 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A1 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A2 = CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D5 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A4 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C2 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A5 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B1 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B2 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C5 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A3 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A4 = CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A5 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A6 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C1 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B2 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B4 = CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B5 = CLBLM_R_X7Y150_SLICE_X9Y150_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B6 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A1 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A2 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A3 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A6 = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B1 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B2 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B4 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B5 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A1 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A3 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A5 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A6 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_AX = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B1 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B2 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B4 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_A5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C3 = CLBLM_R_X5Y144_SLICE_X6Y144_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C4 = CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D2 = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D3 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C5 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D4 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D2 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D3 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D4 = CLBLM_L_X12Y141_SLICE_X16Y141_C5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D6 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C6 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A2 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A3 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A4 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C5 = CLBLM_R_X11Y151_SLICE_X15Y151_CQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B5 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A2 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A5 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A6 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B2 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B4 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B6 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C1 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C2 = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C5 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D1 = CLBLM_L_X12Y144_SLICE_X16Y144_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D2 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D3 = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D6 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A2 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A3 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A4 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A5 = CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A6 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B1 = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B3 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B5 = CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B6 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C2 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C3 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C4 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D3 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D4 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B5 = CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B6 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C1 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D5 = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D6 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A2 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A4 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A5 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B1 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B2 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B4 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B5 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B6 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C1 = CLBLM_L_X12Y143_SLICE_X16Y143_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C2 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C5 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D2 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D3 = CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D4 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D5 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D6 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X12Y143_SLICE_X16Y143_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A1 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A3 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A4 = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B1 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B2 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B3 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B6 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_BX = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C2 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C4 = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C5 = CLBLM_R_X5Y143_SLICE_X6Y143_B5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D3 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D4 = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D5 = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D6 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A1 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A2 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A3 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A4 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A5 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B1 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B2 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B4 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B6 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C2 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C3 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C5 = CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D1 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D4 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D5 = CLBLM_L_X8Y144_SLICE_X10Y144_DQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A2 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A3 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A4 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A5 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A6 = 1'b1;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B1 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B2 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B5 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C2 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C3 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C5 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C6 = CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C3 = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D1 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D2 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D3 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C6 = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X12Y143_SLICE_X16Y143_C5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A3 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A6 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B2 = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B5 = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B6 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C2 = CLBLM_L_X12Y144_SLICE_X16Y144_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C5 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D2 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A1 = CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A3 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A4 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A6 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_AX = CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B3 = CLBLM_L_X8Y144_SLICE_X10Y144_DQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_CQ;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B5 = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C2 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C3 = CLBLM_L_X8Y141_SLICE_X10Y141_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C4 = CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D1 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D2 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D4 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D5 = CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D2 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C3 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D4 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D5 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C5 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A1 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C1 = CLBLM_R_X11Y141_SLICE_X14Y141_B5Q;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A4 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A5 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A6 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C2 = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B5 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C5 = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A1 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A3 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A4 = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B2 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B3 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B4 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B5 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C1 = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C2 = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C3 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C4 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C5 = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C6 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D6 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A1 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A2 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A4 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D3 = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B2 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B5 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D4 = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B6 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C1 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C2 = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C3 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D6 = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D1 = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D2 = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D3 = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D4 = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D5 = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D6 = CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D6 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X37Y143_SLICE_X56Y143_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C4 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C5 = CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C6 = CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A2 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A3 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A4 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D1 = CLBLM_R_X13Y148_SLICE_X19Y148_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D2 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B1 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B2 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B3 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B4 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B5 = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B6 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C1 = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C2 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C4 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C5 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C6 = CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D1 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D2 = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D3 = CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D4 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D5 = CLBLM_L_X10Y149_SLICE_X12Y149_DQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D6 = CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A1 = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A2 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A3 = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A4 = CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A5 = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A6 = CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B1 = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B2 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B3 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B4 = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B5 = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B6 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_R_X13Y147_SLICE_X18Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C1 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C2 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C3 = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C4 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C5 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C6 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D1 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D3 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D4 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D6 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D2 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D3 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B4 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B5 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B6 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C3 = CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C5 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D5 = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A1 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A2 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A3 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A4 = CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A6 = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B2 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B3 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B5 = CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C2 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C4 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C5 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C6 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D1 = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D2 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D3 = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D4 = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D5 = CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D6 = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A2 = CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A3 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A4 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B2 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B3 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B5 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B6 = CLBLM_R_X7Y143_SLICE_X9Y143_DQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C1 = CLBLM_R_X11Y144_SLICE_X14Y144_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C3 = CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C4 = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C5 = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C6 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D1 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D2 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D3 = CLBLM_L_X8Y148_SLICE_X10Y148_DQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D4 = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D5 = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D6 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D1 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A2 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A4 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A5 = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A6 = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B4 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C1 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C3 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C4 = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C5 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C6 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D1 = CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D3 = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D4 = CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D5 = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D6 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A1 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A2 = CLBLM_R_X11Y147_SLICE_X15Y147_D5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A6 = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B5 = CLBLM_R_X11Y142_SLICE_X14Y142_C5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B1 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B2 = CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B4 = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B5 = CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B6 = CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C2 = CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C3 = CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C4 = CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C5 = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C6 = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D1 = CLBLM_L_X12Y147_SLICE_X17Y147_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D2 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D3 = CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D4 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D5 = CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D6 = CLBLM_R_X5Y150_SLICE_X6Y150_AO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C5 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C6 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D4 = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A4 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B3 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B4 = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B5 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C5 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D5 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B2 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B5 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B6 = CLBLM_R_X7Y150_SLICE_X9Y150_BQ;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C4 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C5 = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C6 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D1 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D4 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D5 = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D6 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D6 = CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C6 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C3 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C4 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C5 = CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C6 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B5 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C4 = CLBLM_L_X12Y152_SLICE_X17Y152_CO5;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C5 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B5 = CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C2 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C4 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C5 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C6 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D1 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D2 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D3 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D4 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D5 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C3 = CLBLM_L_X12Y146_SLICE_X17Y146_CQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D6 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_B5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C2 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C3 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C4 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C5 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_R_X13Y151_SLICE_X19Y151_AO5;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A2 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A4 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A5 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B1 = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B3 = CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B4 = CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B5 = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B6 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C2 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C4 = CLBLM_R_X7Y141_SLICE_X9Y141_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C5 = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C6 = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D3 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D4 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D5 = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D6 = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A2 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A4 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A5 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B2 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C2 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B2 = CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D2 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B6 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A3 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A5 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A6 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_AX = CLBLM_R_X3Y144_SLICE_X3Y144_AO5;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_DQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B5 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B6 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C2 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C2 = CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C3 = CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D2 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A1 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A3 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A4 = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A6 = CLBLM_L_X12Y148_SLICE_X17Y148_DQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C6 = CLBLM_L_X12Y141_SLICE_X16Y141_BO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B1 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B2 = CLBLM_L_X12Y139_SLICE_X17Y139_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_B5Q;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C1 = CLBLM_L_X12Y141_SLICE_X17Y141_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C2 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C4 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_A1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A3 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_A2 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_A3 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_A4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A4 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D1 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D2 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D3 = CLBLM_L_X12Y139_SLICE_X17Y139_DQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_B1 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_B2 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_B3 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_B4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A1 = CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A2 = CLBLM_L_X12Y141_SLICE_X16Y141_CQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A3 = CLBLM_L_X12Y139_SLICE_X16Y139_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A4 = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A5 = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_C1 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_C2 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_C3 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_C4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B1 = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B2 = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B3 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B5 = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B6 = CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_D1 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_D2 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_D3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C1 = CLBLM_R_X11Y138_SLICE_X14Y138_DO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C2 = CLBLM_L_X12Y141_SLICE_X16Y141_CQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C2 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C4 = CLBLM_L_X12Y139_SLICE_X16Y139_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B2 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C5 = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C6 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_A1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B3 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_A3 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B4 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D1 = CLBLM_R_X11Y138_SLICE_X14Y138_DO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D2 = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D4 = CLBLM_L_X12Y141_SLICE_X16Y141_CQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B5 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B6 = CLBLM_L_X10Y141_SLICE_X12Y141_A5Q;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_C3 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_D1 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_D2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_D3 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_D4 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_D5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C2 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C4 = CLBLM_L_X12Y148_SLICE_X17Y148_DQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C5 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_BQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D3 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D4 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X11Y142_SLICE_X14Y142_C5Q;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A1 = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A3 = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A4 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A5 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A6 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_R_X13Y151_SLICE_X19Y151_AO5;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B1 = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B2 = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B3 = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B4 = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B5 = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C1 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C2 = CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C3 = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C4 = CLBLM_R_X7Y141_SLICE_X9Y141_CQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C6 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D1 = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D2 = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A2 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B2 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B5 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C1 = CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C2 = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C4 = CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C6 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A3 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A4 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A5 = CLBLM_L_X12Y142_SLICE_X17Y142_DQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B2 = CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B3 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B4 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B6 = CLBLM_L_X12Y141_SLICE_X17Y141_BQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C2 = CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C4 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C5 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C6 = CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D1 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D2 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D3 = CLBLM_R_X11Y141_SLICE_X14Y141_B5Q;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D4 = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D6 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A1 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A3 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A4 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A5 = CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B1 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B2 = CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B3 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B4 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B6 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C1 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C2 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C4 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C5 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D1 = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D2 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D4 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D5 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D6 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D1 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A6 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C6 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D6 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A2 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A3 = CLBLM_R_X15Y144_SLICE_X20Y144_AQ;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B6 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C6 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A1 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A2 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A3 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A4 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B1 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B2 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B3 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B4 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C1 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C2 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C3 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C4 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D1 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D2 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D3 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D4 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A4 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C4 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D2 = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D4 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D6 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C5 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A1 = CLBLM_L_X12Y141_SLICE_X17Y141_CQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A3 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A4 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A5 = CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B2 = CLBLM_L_X12Y141_SLICE_X17Y141_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B3 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C2 = CLBLM_L_X12Y141_SLICE_X17Y141_CQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C3 = CLBLM_L_X12Y139_SLICE_X17Y139_DQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C4 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C5 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D1 = CLBLM_L_X12Y139_SLICE_X17Y139_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D2 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D3 = CLBLM_R_X13Y141_SLICE_X18Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D4 = CLBLM_L_X12Y141_SLICE_X17Y141_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D5 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D6 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A2 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A3 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A4 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A5 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D2 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_AX = CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B2 = CLBLM_L_X12Y139_SLICE_X17Y139_BQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B5 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C1 = CLBLM_L_X12Y139_SLICE_X16Y139_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C4 = CLBLM_L_X12Y142_SLICE_X16Y142_A5Q;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C5 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D1 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D2 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D3 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D4 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D6 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B4 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X7Y142_SLICE_X9Y142_B5Q;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B5 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A1 = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A2 = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A3 = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A5 = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A6 = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B2 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C4 = CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C1 = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C2 = CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C3 = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C4 = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C5 = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C6 = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C5 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C6 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D1 = CLBLM_R_X5Y144_SLICE_X7Y144_DQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D2 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D4 = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D5 = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D6 = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A2 = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A3 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A4 = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A5 = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A6 = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B2 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B4 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B6 = CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C1 = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C2 = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C4 = CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C5 = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C6 = CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D1 = CLBLM_R_X5Y143_SLICE_X6Y143_B5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D2 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A1 = CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A3 = CLBLM_L_X12Y142_SLICE_X16Y142_A5Q;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C3 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B4 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B5 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C1 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C2 = CLBLM_L_X12Y142_SLICE_X17Y142_CQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C3 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D1 = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D2 = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D3 = CLBLM_L_X12Y142_SLICE_X17Y142_DQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B3 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A3 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A4 = CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A5 = CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_AX = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B1 = CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B2 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B3 = CLBLM_L_X12Y144_SLICE_X16Y144_DQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B4 = CLBLM_R_X11Y142_SLICE_X14Y142_B5Q;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D1 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D2 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D3 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C2 = CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C3 = CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C5 = CLBLM_R_X13Y145_SLICE_X18Y145_AQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C6 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D4 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D1 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D2 = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D3 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D5 = CLBLM_L_X12Y147_SLICE_X16Y147_DQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D6 = CLBLM_R_X13Y142_SLICE_X18Y142_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D3 = CLBLM_L_X10Y149_SLICE_X12Y149_DQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D2 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D3 = CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B1 = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B2 = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B3 = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B4 = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B5 = CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C1 = CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C2 = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C4 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C5 = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A1 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D2 = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D3 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D4 = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D5 = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D6 = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A4 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B2 = CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B3 = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B4 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B5 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B6 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C2 = CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C4 = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B2 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D2 = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D3 = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D4 = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D5 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A3 = CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A5 = CLBLM_R_X13Y142_SLICE_X18Y142_CQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B2 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B4 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B5 = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C2 = CLBLM_L_X12Y148_SLICE_X17Y148_CQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C5 = CLBLM_L_X8Y143_SLICE_X11Y143_C5Q;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D3 = CLBLM_L_X12Y143_SLICE_X16Y143_B5Q;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D5 = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D6 = CLBLM_L_X12Y143_SLICE_X17Y143_DQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A3 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A5 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_CQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B1 = CLBLM_L_X12Y143_SLICE_X17Y143_A5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B3 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B4 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C1 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C4 = CLBLM_R_X13Y145_SLICE_X18Y145_BQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C5 = CLBLM_L_X12Y143_SLICE_X16Y143_B5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D2 = CLBLM_L_X12Y143_SLICE_X17Y143_A5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D3 = CLBLM_L_X12Y144_SLICE_X16Y144_DQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D4 = CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D6 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D1 = 1'b1;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A2 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B1 = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B3 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C2 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C3 = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C4 = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C5 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C6 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D2 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D3 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D4 = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D5 = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D6 = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_R_X13Y147_SLICE_X18Y147_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B4 = CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B5 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B6 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B1 = CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B2 = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B3 = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B4 = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B5 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C6 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_A5 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_A6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D2 = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D3 = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D4 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D5 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D6 = CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A1 = CLBLM_R_X13Y145_SLICE_X18Y145_BQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A3 = CLBLM_R_X13Y145_SLICE_X18Y145_CQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A4 = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A5 = CLBLM_R_X13Y145_SLICE_X19Y145_CQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_AX = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B1 = CLBLM_L_X12Y144_SLICE_X17Y144_BQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B4 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B6 = CLBLM_L_X12Y146_SLICE_X17Y146_BQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C1 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C2 = CLBLM_L_X12Y144_SLICE_X17Y144_CQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C4 = CLBLM_L_X12Y144_SLICE_X17Y144_BQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_B5 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D1 = CLBLM_R_X13Y143_SLICE_X19Y143_BQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D2 = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D3 = CLBLM_R_X13Y146_SLICE_X19Y146_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D4 = CLBLM_R_X13Y145_SLICE_X18Y145_DQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D5 = CLBLM_L_X12Y145_SLICE_X17Y145_DQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D6 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A2 = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A3 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A5 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_AX = CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B1 = CLBLM_R_X13Y145_SLICE_X18Y145_DQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B2 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B3 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B6 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C3 = CLBLM_R_X13Y141_SLICE_X18Y141_A5Q;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C4 = CLBLM_L_X12Y145_SLICE_X17Y145_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C5 = CLBLM_L_X8Y143_SLICE_X11Y143_C5Q;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C6 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_C5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_C6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D2 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D6 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_D4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_D5 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X57Y143_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_A5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_A6 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B3 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B4 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C3 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C4 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C5 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_B1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D3 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D4 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D6 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_B2 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_B3 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_B4 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A6 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_B5 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_B6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B5 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C3 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C4 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D3 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D4 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D6 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_C1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A3 = CLBLM_L_X12Y145_SLICE_X17Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A6 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_C2 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B2 = CLBLM_L_X12Y145_SLICE_X17Y145_BQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B3 = CLBLM_L_X12Y145_SLICE_X17Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B4 = CLBLM_L_X12Y147_SLICE_X17Y147_BQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_C5 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C2 = CLBLM_L_X12Y145_SLICE_X17Y145_CQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C3 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C6 = CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_C6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D2 = CLBLM_R_X13Y145_SLICE_X18Y145_BQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D3 = CLBLM_L_X12Y145_SLICE_X17Y145_DQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A2 = CLBLM_R_X13Y145_SLICE_X18Y145_DQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A3 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A4 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A6 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B1 = CLBLM_L_X12Y143_SLICE_X17Y143_B5Q;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B2 = CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B4 = CLBLM_L_X12Y145_SLICE_X16Y145_CQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C2 = CLBLM_L_X12Y145_SLICE_X16Y145_CQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C3 = CLBLM_L_X12Y139_SLICE_X16Y139_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C4 = CLBLM_R_X11Y145_SLICE_X15Y145_DQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D3 = CLBLM_L_X12Y147_SLICE_X16Y147_DQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D4 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D5 = CLBLM_R_X11Y145_SLICE_X15Y145_CQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D6 = 1'b1;
  assign CLBLM_R_X37Y143_SLICE_X56Y143_D6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C1 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C2 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C6 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D1 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D6 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A1 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A3 = CLBLM_L_X12Y146_SLICE_X17Y146_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A5 = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B2 = CLBLM_L_X12Y146_SLICE_X17Y146_BQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B5 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_DQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C2 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C4 = CLBLM_L_X12Y146_SLICE_X17Y146_BQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D3 = CLBLM_R_X13Y146_SLICE_X19Y146_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D4 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A1 = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A4 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A6 = CLBLM_L_X12Y144_SLICE_X16Y144_A5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_AX = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B2 = CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B5 = CLBLM_L_X12Y144_SLICE_X16Y144_CO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B6 = CLBLM_L_X12Y146_SLICE_X16Y146_A5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C1 = CLBLM_R_X13Y145_SLICE_X18Y145_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C4 = CLBLM_R_X13Y145_SLICE_X18Y145_CQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D2 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D3 = CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D6 = CLBLM_L_X12Y145_SLICE_X16Y145_DO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C6 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y135_SLICE_X0Y135_AO5;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y135_SLICE_X0Y135_BO5;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A6 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D6 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A1 = CLBLM_L_X12Y143_SLICE_X17Y143_DQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A3 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A6 = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C3 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D1 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A2 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D3 = CLBLM_L_X12Y146_SLICE_X17Y146_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D4 = CLBLM_L_X12Y143_SLICE_X17Y143_DQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_DQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A3 = CLBLM_L_X12Y147_SLICE_X17Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A4 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B1 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B2 = CLBLM_L_X12Y147_SLICE_X17Y147_BQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B3 = CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B2 = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A1 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C6 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C2 = CLBLM_L_X12Y147_SLICE_X17Y147_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D2 = CLBLM_L_X12Y147_SLICE_X17Y147_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A3 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A4 = CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A5 = CLBLM_R_X13Y148_SLICE_X18Y148_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B1 = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B2 = CLBLM_L_X12Y147_SLICE_X16Y147_BQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A2 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A4 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A6 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C2 = CLBLM_L_X12Y147_SLICE_X16Y147_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B2 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B5 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D4 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B6 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B6 = 1'b1;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D3 = CLBLM_L_X10Y149_SLICE_X13Y149_DQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C3 = CLBLM_L_X12Y149_SLICE_X16Y149_DQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A1 = CLBLM_R_X11Y141_SLICE_X14Y141_B5Q;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A3 = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A5 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B3 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C6 = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B6 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C3 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C5 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A3 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A5 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D3 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D5 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A6 = CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A3 = CLBLM_R_X13Y141_SLICE_X18Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A5 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_AX = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C3 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B2 = CLBLM_R_X13Y141_SLICE_X18Y141_A5Q;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B4 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B5 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C3 = CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A6 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D3 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D5 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B1 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B2 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A5 = CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A6 = CLBLM_R_X13Y151_SLICE_X18Y151_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C2 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C3 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B2 = CLBLM_R_X13Y147_SLICE_X18Y147_CQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B3 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B5 = CLBLM_L_X12Y148_SLICE_X17Y148_BQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B6 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A1 = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A2 = CLBLM_L_X10Y141_SLICE_X12Y141_A5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A3 = CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A4 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A5 = CLBLM_R_X13Y142_SLICE_X18Y142_A5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A6 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C2 = CLBLM_L_X12Y148_SLICE_X17Y148_CQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B1 = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B2 = CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B3 = CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B4 = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B5 = CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B6 = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D3 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C1 = CLBLM_R_X11Y142_SLICE_X14Y142_CQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C2 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C3 = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C5 = CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C6 = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D5 = CLBLM_R_X13Y148_SLICE_X18Y148_AQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A1 = CLBLM_R_X15Y144_SLICE_X20Y144_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A3 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A4 = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A5 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_AX = CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B1 = CLBLM_L_X12Y149_SLICE_X16Y149_DQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B3 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B4 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B5 = CLBLM_L_X12Y149_SLICE_X17Y149_DQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A1 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A3 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A6 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_BX = CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C1 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C3 = CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B3 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B6 = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C1 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C3 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C4 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C5 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_SR = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D4 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D5 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A1 = CLBLM_R_X13Y142_SLICE_X18Y142_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A1 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A3 = CLBLM_R_X13Y146_SLICE_X18Y146_CQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A5 = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_AX = CLBLM_R_X13Y147_SLICE_X18Y147_DO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B1 = CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B6 = CLBLM_R_X13Y141_SLICE_X18Y141_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C4 = CLBLM_R_X13Y142_SLICE_X18Y142_A5Q;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A2 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A4 = CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C5 = CLBLM_L_X12Y144_SLICE_X16Y144_DQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D1 = CLBLM_R_X13Y146_SLICE_X18Y146_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D2 = CLBLM_R_X13Y142_SLICE_X18Y142_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D3 = CLBLM_L_X12Y148_SLICE_X17Y148_CQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D5 = CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D6 = CLBLM_R_X13Y143_SLICE_X19Y143_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A3 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B1 = CLBLM_L_X12Y145_SLICE_X16Y145_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B3 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B6 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A3 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A4 = CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A5 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A6 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B1 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B2 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B4 = CLBLM_L_X12Y149_SLICE_X17Y149_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B5 = CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B6 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C4 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A1 = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A2 = CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A3 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A4 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A5 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A6 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C1 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C2 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B1 = CLBLM_R_X11Y141_SLICE_X14Y141_B5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B3 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B4 = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B5 = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B6 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C1 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C2 = CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C3 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C4 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C6 = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D5 = CLBLM_L_X12Y148_SLICE_X17Y148_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A1 = CLBLM_L_X10Y149_SLICE_X12Y149_DQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A2 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A3 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A4 = CLBLM_L_X12Y150_SLICE_X17Y150_CQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A6 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D2 = CLBLM_L_X10Y141_SLICE_X12Y141_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D3 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D4 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D6 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B1 = CLBLM_L_X12Y146_SLICE_X17Y146_CQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B2 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B3 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B5 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A3 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A4 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A6 = CLBLM_L_X12Y139_SLICE_X16Y139_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C1 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B3 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B4 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B5 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B6 = CLBLM_R_X13Y141_SLICE_X18Y141_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D2 = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C2 = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C3 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C4 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C5 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C6 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D3 = CLBLM_L_X12Y149_SLICE_X16Y149_DQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D4 = CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B3 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D1 = CLBLM_R_X11Y139_SLICE_X14Y139_DO5;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D2 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D3 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_C5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D6 = CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B1 = CLBLM_L_X10Y143_SLICE_X13Y143_DQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B2 = CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C1 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C2 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A2 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A6 = CLBLM_R_X13Y143_SLICE_X19Y143_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B2 = CLBLM_R_X13Y143_SLICE_X19Y143_BQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B4 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B5 = CLBLM_R_X13Y146_SLICE_X18Y146_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B6 = CLBLM_R_X13Y143_SLICE_X19Y143_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C2 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C4 = CLBLM_L_X12Y145_SLICE_X17Y145_BQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C5 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C6 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D1 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D2 = CLBLM_R_X13Y145_SLICE_X19Y145_BQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D3 = CLBLM_R_X13Y145_SLICE_X19Y145_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D4 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D5 = CLBLM_R_X13Y143_SLICE_X19Y143_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D6 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C5 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A3 = CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A6 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B1 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B2 = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B6 = CLBLM_R_X13Y145_SLICE_X19Y145_CQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C1 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C2 = CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C4 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D2 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C5 = CLBLM_L_X12Y145_SLICE_X17Y145_CQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C6 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D3 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D1 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D2 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D3 = CLBLM_L_X12Y145_SLICE_X17Y145_CQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D4 = CLBLM_R_X13Y145_SLICE_X19Y145_CQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D5 = CLBLM_R_X13Y145_SLICE_X19Y145_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D6 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A1 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A1 = CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A2 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A3 = CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A4 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A6 = CLBLM_L_X12Y151_SLICE_X17Y151_AO5;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B2 = CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B4 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B5 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B6 = CLBLM_L_X12Y150_SLICE_X17Y150_DQ;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A1 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A4 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A5 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C2 = CLBLM_L_X12Y150_SLICE_X17Y150_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B1 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B5 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D3 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D4 = CLBLM_L_X12Y150_SLICE_X17Y150_DQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C2 = CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C3 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C5 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D5 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D6 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A1 = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A2 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A5 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D1 = CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D2 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D3 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D4 = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D5 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_AX = CLBLM_R_X13Y150_SLICE_X18Y150_AO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B1 = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B4 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A1 = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_BX = CLBLM_R_X13Y151_SLICE_X19Y151_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C1 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C2 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C3 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B1 = CLBLM_L_X10Y140_SLICE_X12Y140_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B4 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B5 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_BX = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D3 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C1 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C2 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C4 = CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C5 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C6 = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D4 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D5 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D6 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D3 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D4 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D5 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D6 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D5 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A1 = CLBLM_R_X13Y145_SLICE_X18Y145_DQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A2 = CLBLM_R_X13Y143_SLICE_X18Y143_DO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A4 = CLBLM_R_X13Y145_SLICE_X18Y145_CQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A5 = CLBLM_R_X13Y146_SLICE_X18Y146_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A6 = CLBLM_L_X12Y148_SLICE_X17Y148_CQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B1 = CLBLM_R_X13Y144_SLICE_X19Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B3 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B4 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B5 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B6 = CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D6 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C2 = CLBLM_L_X12Y145_SLICE_X17Y145_BQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C4 = CLBLM_R_X13Y145_SLICE_X19Y145_BQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C6 = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D1 = CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D4 = CLBLM_R_X13Y146_SLICE_X19Y146_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D6 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A1 = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A2 = CLBLM_R_X13Y144_SLICE_X19Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A3 = CLBLM_R_X13Y144_SLICE_X19Y144_AO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A4 = CLBLM_R_X13Y144_SLICE_X18Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A5 = CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A6 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B1 = CLBLM_R_X13Y143_SLICE_X19Y143_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B2 = CLBLM_R_X13Y145_SLICE_X18Y145_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B3 = CLBLM_R_X13Y145_SLICE_X18Y145_CQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B4 = CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B5 = CLBLM_R_X13Y145_SLICE_X19Y145_CQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B6 = CLBLM_L_X12Y146_SLICE_X17Y146_BQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C1 = CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C2 = CLBLM_L_X12Y146_SLICE_X17Y146_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C4 = CLBLM_L_X12Y144_SLICE_X17Y144_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C5 = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C6 = CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D1 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D2 = CLBLM_L_X12Y144_SLICE_X17Y144_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D3 = CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D4 = CLBLM_L_X12Y146_SLICE_X17Y146_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D5 = CLBLM_R_X13Y143_SLICE_X19Y143_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D6 = CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A1 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A2 = CLBLM_L_X12Y152_SLICE_X16Y152_DO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A3 = CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A4 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A5 = CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_AX = CLBLM_L_X12Y150_SLICE_X17Y150_DQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B1 = CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B2 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B3 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B4 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B5 = CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B6 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A1 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C4 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C5 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C6 = CLBLM_L_X12Y150_SLICE_X17Y150_DQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A4 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A5 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B3 = CLBLM_R_X13Y143_SLICE_X19Y143_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B5 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B6 = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D5 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D6 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D1 = CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C1 = CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C2 = CLBLM_L_X10Y141_SLICE_X12Y141_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C4 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C5 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C6 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A2 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A5 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D1 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D3 = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D4 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D6 = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B5 = CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B6 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_AX = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B1 = CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B2 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B3 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B4 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_B5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C4 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C5 = CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C6 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A3 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C2 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_AX = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B3 = CLBLM_L_X10Y149_SLICE_X13Y149_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B4 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B5 = CLBLM_L_X12Y142_SLICE_X17Y142_DQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CX = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D5 = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D1 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C2 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C4 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C5 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_SR = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D2 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D4 = CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D6 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A4 = CLBLM_R_X11Y149_SLICE_X14Y149_A5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A3 = CLBLM_R_X13Y145_SLICE_X19Y145_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A4 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A6 = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B2 = CLBLM_R_X13Y145_SLICE_X19Y145_BQ;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B3 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B6 = CLBLM_R_X13Y145_SLICE_X18Y145_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C2 = CLBLM_R_X13Y145_SLICE_X19Y145_CQ;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C3 = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C6 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A6 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D1 = CLBLM_R_X11Y145_SLICE_X15Y145_DQ;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D4 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D6 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A3 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A2 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A3 = CLBLM_R_X13Y145_SLICE_X18Y145_AQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A5 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B1 = CLBLM_R_X13Y143_SLICE_X19Y143_BQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B2 = CLBLM_R_X13Y145_SLICE_X18Y145_BQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B4 = CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C2 = CLBLM_R_X13Y145_SLICE_X18Y145_CQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C4 = CLBLM_R_X13Y146_SLICE_X19Y146_AQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C5 = CLBLM_L_X12Y148_SLICE_X17Y148_DQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C4 = CLBLM_L_X12Y150_SLICE_X17Y150_CQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D1 = CLBLM_R_X13Y145_SLICE_X19Y145_AQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D3 = CLBLM_R_X13Y145_SLICE_X18Y145_DQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C6 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B3 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A1 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A2 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A3 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A4 = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A6 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B1 = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B2 = CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B4 = CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D1 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D2 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D6 = 1'b1;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A1 = CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A2 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A3 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A4 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B1 = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B2 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B3 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B4 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B6 = CLBLM_L_X10Y149_SLICE_X13Y149_CQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C1 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C2 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C3 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C5 = CLBLM_R_X13Y152_SLICE_X18Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A1 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A2 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D1 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D2 = CLBLM_L_X12Y150_SLICE_X17Y150_CQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D3 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D4 = CLBLM_R_X13Y152_SLICE_X18Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D5 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D6 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B4 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_BX = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C2 = CLBLM_R_X13Y142_SLICE_X18Y142_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A1 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A3 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A4 = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A5 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A6 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D1 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B2 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B4 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B5 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B6 = CLBLM_L_X12Y154_SLICE_X16Y154_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D4 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D5 = CLBLM_L_X10Y142_SLICE_X13Y142_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C4 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C5 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A5 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A6 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C2 = CLBLM_L_X12Y152_SLICE_X17Y152_CO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B1 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B2 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D2 = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D3 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B6 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D5 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D1 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C2 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C4 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C6 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D1 = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D2 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D5 = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A1 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A3 = CLBLM_R_X13Y146_SLICE_X19Y146_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A4 = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C4 = CLBLM_R_X13Y147_SLICE_X18Y147_CQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C6 = CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A2 = CLBLM_L_X12Y144_SLICE_X17Y144_CQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A3 = CLBLM_R_X13Y146_SLICE_X18Y146_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A4 = CLBLM_R_X13Y147_SLICE_X18Y147_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B1 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B3 = CLBLL_L_X4Y140_SLICE_X4Y140_BQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B5 = CLBLM_R_X13Y146_SLICE_X18Y146_CQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C2 = CLBLM_R_X13Y146_SLICE_X18Y146_CQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C5 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D1 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A1 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A3 = CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A4 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A5 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_AX = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B2 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B3 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B4 = CLBLL_L_X4Y139_SLICE_X4Y139_DO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B5 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B6 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C2 = CLBLL_L_X4Y139_SLICE_X5Y139_AO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C3 = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C5 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C6 = CLBLM_L_X8Y142_SLICE_X11Y142_A5Q;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B3 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D4 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D3 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A1 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A2 = CLBLM_L_X12Y146_SLICE_X17Y146_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A4 = CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A5 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B1 = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B2 = CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B3 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B4 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B5 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B6 = CLBLM_R_X13Y152_SLICE_X18Y152_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A1 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A2 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A3 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C1 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C2 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C3 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C4 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C5 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C6 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B1 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B2 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B3 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B5 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D1 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C1 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C2 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C2 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C6 = CLBLM_L_X10Y143_SLICE_X13Y143_CQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D1 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D2 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A4 = CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A5 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D4 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D2 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B3 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B4 = CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B5 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B6 = CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D3 = CLBLM_L_X10Y142_SLICE_X13Y142_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A2 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C3 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C4 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C5 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C6 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A3 = CLBLM_R_X5Y143_SLICE_X6Y143_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A4 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B1 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B4 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B5 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D1 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D5 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D6 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C5 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D3 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D4 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D1 = CLBLM_L_X12Y141_SLICE_X16Y141_BO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D2 = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D5 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D6 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D6 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A2 = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A4 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A2 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A3 = CLBLM_R_X13Y147_SLICE_X18Y147_AQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A5 = CLBLM_L_X12Y147_SLICE_X16Y147_BQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B1 = CLBLM_R_X13Y148_SLICE_X18Y148_CQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B2 = CLBLM_R_X13Y147_SLICE_X18Y147_BQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B4 = CLBLM_R_X13Y147_SLICE_X18Y147_DO5;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B6 = CLBLM_L_X12Y144_SLICE_X17Y144_CQ;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C4 = CLBLM_R_X13Y146_SLICE_X18Y146_BO5;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C5 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C6 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D2 = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D3 = CLBLM_R_X13Y148_SLICE_X18Y148_BQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D4 = CLBLM_L_X12Y146_SLICE_X16Y146_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A5 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D5 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A6 = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A1 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A2 = CLBLL_L_X4Y139_SLICE_X4Y139_DO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A3 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A4 = CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A6 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C2 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_AX = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B1 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B2 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B3 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B4 = CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B5 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C2 = CLBLL_L_X4Y140_SLICE_X4Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C3 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C5 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C6 = CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D1 = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D2 = CLBLL_L_X4Y139_SLICE_X5Y139_AO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A2 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A3 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A4 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A5 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A6 = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A3 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B4 = CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B5 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C1 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C2 = CLBLM_L_X10Y142_SLICE_X13Y142_B5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C3 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C4 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C5 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D1 = CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D4 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D5 = CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D6 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B1 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B2 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B3 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B4 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A2 = CLBLM_R_X11Y142_SLICE_X14Y142_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A3 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A4 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C2 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_B5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B4 = CLBLM_L_X12Y143_SLICE_X17Y143_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C2 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C3 = CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C4 = CLBLM_R_X13Y141_SLICE_X18Y141_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C6 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D3 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D4 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D1 = CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D2 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D4 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D5 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D6 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B1 = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B3 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B4 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_AX = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B4 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A1 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A4 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A6 = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C3 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B3 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B4 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B5 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C1 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C2 = CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C3 = CLBLM_R_X11Y138_SLICE_X14Y138_BO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C4 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C2 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C5 = CLBLM_R_X11Y138_SLICE_X15Y138_BO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C6 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A1 = CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C3 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C4 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D1 = CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D2 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D3 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D4 = CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C5 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D5 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D6 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_AX = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B1 = CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B2 = CLBLM_R_X13Y148_SLICE_X18Y148_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A1 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A5 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C2 = CLBLM_R_X13Y148_SLICE_X18Y148_CQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C3 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B1 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B3 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B4 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B5 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A5 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C2 = CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C4 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C5 = CLBLM_R_X11Y141_SLICE_X14Y141_A5Q;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C6 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D5 = CLBLM_R_X13Y147_SLICE_X18Y147_BQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A1 = CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A2 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A3 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A5 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D1 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B1 = CLBLM_R_X7Y141_SLICE_X8Y141_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B2 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B5 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B6 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D3 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D5 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C1 = CLBLM_L_X8Y146_SLICE_X10Y146_D5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C2 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C4 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C5 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D3 = CLBLM_L_X8Y149_SLICE_X10Y149_DQ;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A1 = CLBLM_R_X5Y141_SLICE_X7Y141_B5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A2 = CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A3 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A4 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A2 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B3 = CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A3 = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B4 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B5 = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B6 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A4 = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A1 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A2 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A4 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A5 = CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A6 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B1 = CLBLM_L_X8Y146_SLICE_X10Y146_DQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B2 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B3 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B4 = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C1 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C2 = CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C6 = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D3 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D1 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D2 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D5 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A4 = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A5 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A6 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B2 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B4 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A4 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C2 = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C3 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C5 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C3 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D3 = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D1 = CLBLM_L_X10Y145_SLICE_X13Y145_B5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D6 = CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X11Y142_SLICE_X14Y142_C5Q;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X4Y140_SLICE_X4Y140_BQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A1 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A2 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A3 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A6 = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C3 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B2 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B4 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B5 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D2 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C1 = CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C2 = CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C3 = CLBLM_L_X8Y141_SLICE_X10Y141_C5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C4 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C5 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C6 = CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D4 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A1 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A2 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A3 = CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A4 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A5 = CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D1 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D2 = CLBLM_L_X12Y139_SLICE_X17Y139_DQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D5 = CLBLM_L_X12Y141_SLICE_X17Y141_CQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D6 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B1 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B2 = CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B3 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B4 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A1 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A4 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A5 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C3 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B1 = CLBLM_L_X12Y148_SLICE_X17Y148_DQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B3 = CLBLM_L_X12Y139_SLICE_X16Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B5 = CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D2 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C2 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C3 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C4 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C5 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A1 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A3 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A5 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B1 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B2 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B3 = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B4 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D2 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D3 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C1 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C2 = CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C5 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C6 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D2 = CLBLM_R_X5Y143_SLICE_X6Y143_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D4 = CLBLM_L_X8Y146_SLICE_X10Y146_D5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D5 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D6 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A1 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A2 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A4 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A5 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B1 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B2 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B3 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B4 = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B5 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B6 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C1 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C2 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C3 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C4 = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C5 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A1 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A2 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A4 = CLBLM_R_X11Y142_SLICE_X14Y142_B5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A5 = CLBLM_L_X10Y149_SLICE_X13Y149_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A6 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B1 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D2 = CLBLM_R_X13Y142_SLICE_X18Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D5 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D6 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B2 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B4 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B5 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B6 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C1 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C2 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C3 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C4 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C5 = CLBLM_R_X15Y144_SLICE_X20Y144_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C6 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D1 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D2 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D3 = CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D4 = CLBLM_L_X12Y146_SLICE_X17Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D5 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D6 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A3 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A4 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A6 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B1 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B2 = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B6 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C1 = CLBLM_R_X13Y142_SLICE_X18Y142_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C3 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C4 = CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D1 = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D3 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D4 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D6 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A2 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A3 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B2 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B3 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A1 = CLBLM_L_X12Y141_SLICE_X16Y141_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A2 = CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A3 = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A4 = CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A5 = CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C2 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C3 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B1 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B3 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B4 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B5 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B6 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D2 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C1 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C2 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C3 = CLBLM_R_X11Y142_SLICE_X14Y142_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C4 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C5 = CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C6 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D3 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A4 = CLBLM_R_X13Y148_SLICE_X18Y148_A5Q;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D2 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D3 = CLBLM_R_X13Y142_SLICE_X18Y142_A5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D4 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D5 = CLBLM_L_X8Y141_SLICE_X10Y141_C5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B2 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A1 = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A2 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A3 = CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A4 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C2 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C3 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B2 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C3 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B6 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C4 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A2 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A3 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A4 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A5 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A6 = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_AX = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C6 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B2 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B3 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B5 = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D1 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C1 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C2 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C3 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C5 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D3 = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D4 = CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D5 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D6 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D1 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D2 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D4 = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D6 = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A1 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A2 = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A3 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A5 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A6 = CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B1 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B3 = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B4 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B5 = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B6 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_DQ;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C1 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C4 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C5 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C6 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A1 = CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A2 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A3 = CLBLM_R_X15Y144_SLICE_X20Y144_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A4 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A5 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D2 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D4 = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D6 = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A6 = CLBLM_R_X11Y142_SLICE_X14Y142_B5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B1 = CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B3 = CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B4 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B5 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B6 = CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C1 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C3 = CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C4 = CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C6 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A5 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A5 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D1 = CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D2 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D3 = CLBLM_R_X11Y151_SLICE_X15Y151_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D4 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D5 = CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D6 = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A2 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A3 = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A4 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A6 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B2 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B5 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C3 = CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C1 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B3 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C2 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D1 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D2 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D3 = CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B6 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A2 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A4 = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B1 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B2 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B3 = CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B4 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B5 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B6 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A2 = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A3 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A4 = CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C1 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C2 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B2 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B3 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B4 = CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B5 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C2 = CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C3 = CLBLM_R_X13Y142_SLICE_X18Y142_A5Q;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C4 = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C5 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C6 = CLBLM_R_X13Y141_SLICE_X18Y141_A5Q;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D4 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A2 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A3 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D3 = CLBLM_R_X11Y142_SLICE_X14Y142_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D4 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D5 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D6 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A6 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B1 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B2 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B3 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A2 = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A3 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A6 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D4 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_AX = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C1 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B1 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B4 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B5 = CLBLM_R_X11Y141_SLICE_X14Y141_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A3 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A4 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B1 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B2 = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B3 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B4 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B5 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B6 = CLBLM_L_X8Y144_SLICE_X10Y144_DQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C4 = CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D2 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D3 = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D4 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D5 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A1 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A2 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A3 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A5 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A6 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B2 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B5 = CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B6 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C1 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C2 = CLBLM_L_X8Y144_SLICE_X10Y144_DQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C3 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C4 = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C5 = CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D3 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D4 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D5 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D6 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A2 = CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A3 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A5 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B1 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B2 = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B3 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B4 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B5 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B6 = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C1 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C2 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C3 = CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C4 = CLBLM_R_X11Y149_SLICE_X14Y149_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C5 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C6 = CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D1 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D2 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D6 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A1 = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A2 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A6 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B1 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B2 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B4 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B5 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B6 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C2 = CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C3 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C5 = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C6 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D4 = CLBLM_R_X11Y149_SLICE_X14Y149_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D6 = CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = CLBLM_R_X13Y147_SLICE_X18Y147_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A4 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B4 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A4 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A5 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A6 = CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C2 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D4 = CLBLM_R_X13Y147_SLICE_X18Y147_CQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B2 = CLBLM_L_X10Y142_SLICE_X13Y142_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B3 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B4 = CLBLM_L_X12Y142_SLICE_X17Y142_CQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D5 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C3 = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C4 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C6 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A2 = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A3 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A4 = CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D1 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D3 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D4 = CLBLM_L_X12Y139_SLICE_X17Y139_DQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A6 = CLBLM_R_X13Y148_SLICE_X18Y148_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B1 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B2 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B3 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A1 = CLBLM_R_X13Y145_SLICE_X19Y145_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A2 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A3 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A4 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A6 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C1 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C2 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C3 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B1 = CLBLM_R_X11Y142_SLICE_X14Y142_B5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A2 = CLBLM_L_X8Y144_SLICE_X10Y144_DQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A3 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A4 = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A6 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B2 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B1 = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B2 = CLBLM_L_X12Y145_SLICE_X17Y145_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B3 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C1 = CLBLM_L_X12Y144_SLICE_X17Y144_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C2 = CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D6 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D2 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D3 = CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D1 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D2 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D4 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C4 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C6 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A3 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A4 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A6 = CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B1 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B2 = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B3 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B4 = CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B5 = CLBLM_L_X12Y141_SLICE_X16Y141_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B6 = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B6 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C1 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C3 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C4 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C5 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C6 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A4 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B3 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B4 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B6 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C3 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C4 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D2 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D5 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A4 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A6 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D3 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D4 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B4 = CLBLM_R_X13Y151_SLICE_X18Y151_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C4 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C6 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A1 = CLBLM_L_X12Y143_SLICE_X17Y143_B5Q;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A3 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A4 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D5 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B3 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B4 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C3 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C4 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A3 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A4 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B5 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B6 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D3 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D4 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C4 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C5 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A2 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B3 = CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B4 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D2 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D5 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C1 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C3 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D1 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D2 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B1 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B2 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B4 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B6 = CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A1 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A2 = CLBLM_L_X8Y143_SLICE_X11Y143_C5Q;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_DQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A4 = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A6 = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C4 = CLBLM_L_X8Y142_SLICE_X11Y142_A5Q;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B2 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B3 = CLBLM_L_X12Y147_SLICE_X16Y147_DQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B4 = CLBLM_L_X12Y143_SLICE_X17Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C5 = CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B5 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B6 = CLBLM_R_X13Y142_SLICE_X18Y142_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C1 = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C3 = CLBLM_L_X10Y149_SLICE_X13Y149_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C6 = CLBLM_L_X10Y142_SLICE_X13Y142_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C2 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D1 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D2 = CLBLM_R_X13Y142_SLICE_X18Y142_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D4 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C3 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D5 = CLBLM_L_X12Y147_SLICE_X16Y147_DQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D6 = CLBLM_L_X12Y143_SLICE_X17Y143_CQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A2 = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A3 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A6 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A1 = CLBLL_L_X4Y145_SLICE_X4Y145_B5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C6 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B1 = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B2 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B3 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B4 = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B5 = CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B6 = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C5 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D4 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D1 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_A5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D1 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D2 = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D3 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D4 = CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D6 = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D4 = CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D5 = CLBLM_R_X11Y147_SLICE_X15Y147_BQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_A5Q;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D3 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A2 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A3 = CLBLM_R_X5Y145_SLICE_X6Y145_C5Q;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A5 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D5 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B1 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B2 = CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B3 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B4 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B5 = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B6 = CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C1 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C2 = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C5 = CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C6 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D1 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D3 = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D4 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D6 = CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A1 = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A2 = CLBLM_R_X11Y144_SLICE_X14Y144_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A3 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A5 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B1 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B2 = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B3 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B4 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B5 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B6 = CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A3 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C4 = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C5 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C6 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A5 = CLBLM_R_X5Y144_SLICE_X7Y144_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A6 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C1 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C2 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B1 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B2 = CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B4 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D2 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B6 = CLBLM_R_X7Y148_SLICE_X9Y148_D5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D5 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D6 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C1 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C3 = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C4 = CLBLM_R_X7Y148_SLICE_X9Y148_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C5 = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C6 = CLBLM_R_X7Y140_SLICE_X9Y140_AO5;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A2 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A3 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A4 = CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A5 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B5 = CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B6 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D6 = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B1 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B2 = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B3 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C4 = CLBLM_R_X13Y148_SLICE_X19Y148_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C5 = CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A2 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A3 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A4 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A6 = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B2 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D1 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D2 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C2 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C3 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C6 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D5 = CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D1 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D2 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D3 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D5 = CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D6 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A3 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A6 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B1 = CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B4 = CLBLM_R_X11Y144_SLICE_X15Y144_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B5 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C2 = CLBLM_R_X11Y144_SLICE_X15Y144_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C4 = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C6 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D2 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D5 = CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D6 = CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A1 = CLBLM_L_X10Y149_SLICE_X13Y149_CQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A2 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A2 = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A3 = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A4 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A5 = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A6 = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B2 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B6 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B1 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B2 = CLBLM_R_X11Y144_SLICE_X14Y144_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C1 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C4 = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C5 = CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C6 = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C1 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C5 = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D3 = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D4 = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D6 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D1 = CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D3 = CLBLM_L_X12Y141_SLICE_X16Y141_BO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D6 = CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A3 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A4 = CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A5 = CLBLM_R_X5Y144_SLICE_X7Y144_DQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B5 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A3 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A4 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A6 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C1 = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C2 = CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C6 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C3 = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C4 = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C5 = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B4 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C4 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D6 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C6 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D3 = CLBLM_R_X7Y147_SLICE_X9Y147_DQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D4 = CLBLM_L_X8Y147_SLICE_X11Y147_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A1 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A2 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A4 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A5 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B1 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B2 = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B3 = CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B4 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B5 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B6 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X37Y143_SLICE_X56Y143_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A2 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C4 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C5 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C6 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A4 = CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C1 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C2 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_AX = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B1 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B5 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D1 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D2 = CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D3 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D4 = CLBLM_L_X10Y152_SLICE_X13Y152_AO5;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D6 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C4 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C6 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A2 = CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A3 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A4 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A6 = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B2 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B4 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C1 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C3 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C4 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C5 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A6 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_AX = CLBLM_L_X8Y141_SLICE_X10Y141_DO5;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B3 = CLBLM_L_X8Y146_SLICE_X10Y146_D5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B5 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C1 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C2 = CLBLM_L_X8Y141_SLICE_X11Y141_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D2 = CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D4 = CLBLM_L_X12Y148_SLICE_X17Y148_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A2 = CLBLM_R_X13Y145_SLICE_X19Y145_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A3 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A6 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B1 = CLBLM_R_X13Y147_SLICE_X18Y147_CQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B2 = CLBLM_R_X11Y142_SLICE_X15Y142_BO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B6 = CLBLM_R_X11Y142_SLICE_X14Y142_DQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C2 = CLBLM_R_X11Y145_SLICE_X15Y145_CQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C3 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C4 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D1 = CLBLM_R_X5Y145_SLICE_X6Y145_C5Q;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D3 = CLBLM_R_X11Y145_SLICE_X15Y145_DQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D5 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A1 = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A3 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B1 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B2 = CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B4 = CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B5 = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B6 = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A5 = CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C1 = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C2 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C5 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B4 = CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B5 = CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C3 = CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C1 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C2 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C4 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D1 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D3 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D4 = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D5 = CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D6 = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C5 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C6 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D2 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D3 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B1 = CLBLM_L_X8Y148_SLICE_X11Y148_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B2 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B3 = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B5 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B6 = CLBLM_R_X5Y144_SLICE_X6Y144_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C2 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C3 = CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C4 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C5 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C6 = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D1 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D1 = CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D3 = CLBLM_L_X8Y149_SLICE_X10Y149_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D4 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D5 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D6 = CLBLM_L_X12Y148_SLICE_X17Y148_D5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A1 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A2 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A3 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A4 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A5 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B1 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A4 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B2 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B3 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B4 = CLBLM_R_X11Y151_SLICE_X14Y151_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B5 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B6 = CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A1 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C4 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_C5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C1 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_AX = CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B1 = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C3 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D1 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C2 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C4 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C6 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A1 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A2 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A3 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A4 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D1 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D4 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B4 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D5 = CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D6 = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B1 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B2 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B3 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A1 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A2 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A3 = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C1 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C3 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B2 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B5 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D1 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D2 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C6 = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D5 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D2 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D3 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D6 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B5 = CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B6 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C6 = 1'b1;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A2 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A6 = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B1 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B3 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C4 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B5 = CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C3 = CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C6 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C4 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C5 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C6 = CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D1 = CLBLM_L_X12Y147_SLICE_X16Y147_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D2 = CLBLM_L_X12Y147_SLICE_X16Y147_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D3 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A2 = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A4 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A6 = CLBLL_L_X4Y145_SLICE_X4Y145_B5Q;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D5 = CLBLM_L_X10Y149_SLICE_X13Y149_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A1 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B2 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B5 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C1 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C3 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C4 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C5 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B1 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B4 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B5 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D2 = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D3 = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D4 = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D5 = CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D6 = CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C3 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C4 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D2 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D1 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D4 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D5 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A2 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A3 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A4 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B1 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B3 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A6 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B4 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B5 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A2 = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C1 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C3 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C6 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C2 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D4 = CLBLM_L_X12Y148_SLICE_X17Y148_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A1 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A4 = CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A5 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B2 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B3 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B4 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C1 = CLBLM_R_X13Y143_SLICE_X19Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D2 = CLBLM_L_X12Y141_SLICE_X16Y141_A5Q;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D5 = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A5 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B2 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C2 = CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C4 = CLBLM_L_X10Y142_SLICE_X13Y142_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D4 = CLBLM_L_X10Y142_SLICE_X13Y142_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D5 = CLBLM_L_X8Y148_SLICE_X10Y148_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A1 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A2 = CLBLM_L_X12Y147_SLICE_X17Y147_CQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A3 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A6 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B2 = CLBLM_R_X11Y147_SLICE_X15Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B3 = CLBLM_R_X13Y147_SLICE_X18Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B6 = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C2 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C3 = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C6 = CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A2 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D3 = CLBLM_R_X11Y147_SLICE_X15Y147_DQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B2 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A4 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A5 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A6 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C2 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B2 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B5 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D2 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C1 = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C2 = CLBLM_R_X11Y151_SLICE_X15Y151_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C3 = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C4 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C5 = CLBLM_R_X11Y147_SLICE_X15Y147_DQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C6 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D3 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D5 = CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D6 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B1 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B6 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A2 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B2 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B6 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C2 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C6 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D2 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D6 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C5 = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A1 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A6 = CLBLM_R_X7Y144_SLICE_X9Y144_DQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_AX = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B1 = CLBLM_L_X8Y145_SLICE_X10Y145_DQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B2 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C1 = CLBLM_L_X10Y144_SLICE_X12Y144_B5Q;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C4 = CLBLM_L_X10Y145_SLICE_X13Y145_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C5 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D1 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D2 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D4 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A3 = CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A4 = CLBLM_L_X12Y144_SLICE_X16Y144_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B2 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B4 = CLBLM_L_X12Y144_SLICE_X16Y144_DQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B6 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C4 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C6 = CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D2 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D3 = CLBLM_L_X8Y144_SLICE_X10Y144_DQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D6 = CLBLM_L_X10Y144_SLICE_X12Y144_B5Q;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A1 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A2 = CLBLM_R_X11Y144_SLICE_X15Y144_CQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A4 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A5 = CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A6 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_AX = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B2 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B4 = CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B6 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C2 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C3 = CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C4 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D1 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D2 = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D3 = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D5 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D6 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A1 = CLBLM_L_X10Y149_SLICE_X13Y149_DQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A2 = CLBLM_L_X12Y148_SLICE_X17Y148_D5Q;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A5 = CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B1 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B2 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B3 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B4 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C1 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C2 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C3 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C5 = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C6 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D1 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D2 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D3 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D4 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D6 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A1 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A2 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A5 = CLBLM_L_X8Y143_SLICE_X11Y143_C5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B2 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B3 = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A5 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B4 = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B5 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B6 = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C1 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C2 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C3 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C5 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C6 = CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D1 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D3 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D4 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D5 = CLBLM_L_X8Y145_SLICE_X10Y145_DQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D6 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A2 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A3 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A5 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_AX = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
endmodule
