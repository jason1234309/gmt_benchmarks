module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input LIOB33_X0Y123_IOB_X0Y124_IPAD,
  input LIOB33_X0Y125_IOB_X0Y125_IPAD,
  input LIOB33_X0Y125_IOB_X0Y126_IPAD,
  input LIOB33_X0Y127_IOB_X0Y127_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AMUX;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AMUX;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_AMUX;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_BO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_DO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_DO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_AO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_BO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_CO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_DO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_DO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_AO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_BO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_BO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_CO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_CO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_DO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_DO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_BO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_BO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_DO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_DO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffaffffffff)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe00f800f800f000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffb0f0fffff0f0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000777f00000044)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0a000f00)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_DO6),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0c0000ff0f0000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fff0ff50)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I3(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I4(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I5(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3323332340004000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fcf8f0f0)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30003000f500f500)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_CLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(1'b1),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h20202020a0a0f0f0)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_BLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(1'b1),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110010)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_ALUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X2Y116_SLICE_X1Y116_CO6),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff1fff1f1)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_BO6),
.I3(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_DO6),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0abb000000330033)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y121_IOB_X0Y121_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00e000e050405040)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y121_IOB_X0Y121_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000100010000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_DO6),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_BO6),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffffffffffff)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcccecc0f000a00)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020000000a00000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h500000000fffffff)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(1'b1),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffffff7fffff)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fafa0000c8c8)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.I3(1'b1),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I5(RIOB33_X105Y119_IOB_X1Y119_I),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f1ffff)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccc800000005)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffccffafffcc)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(LIOB33_X0Y123_IOB_X0Y123_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(RIOB33_X105Y119_IOB_X1Y120_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h04cc000015dd0000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y121_IOB_X0Y121_I),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110010)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_CO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccdcdcccccccfc)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_DO6),
.I2(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0044c0c4)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfa88facc008800)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y121_IOB_X0Y121_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y119_IOB_X1Y120_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffe8e88080)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cf00aaffbaff)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1100ff003333ff33)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff0011aabb)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0c4c4c4c4c)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(1'b1),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffdcc8f8f8f8f)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccaf8caf8c)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y123_IOB_X0Y123_I),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7fffffffff)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X2Y127_SLICE_X0Y127_AO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010033333333)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_ALUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_DO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_BO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5ffaaaaeeee)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_ALUT (
.I0(CLBLL_L_X2Y127_SLICE_X0Y127_AO6),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_AO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_DO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_CO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_BO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_AO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_DO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_CO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_BO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_ALUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_AO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_DO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_CO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_BO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_AO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000000011111111)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0088008800000008)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y127_IOB_X0Y127_I),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0003055f55575)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c404c5f00400000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcfeffff)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeaeeaaaaaaaa)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_DO6),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafa32fafafa)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c000c000c000d1)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033110000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.I2(1'b1),
.I3(LIOB33_X0Y125_IOB_X0Y126_I),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000c880)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a008a008a008acf)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc000050545050)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff700fffeff00)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044004500)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_CO6),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffaaaaaaa8)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(LIOB33_X0Y121_IOB_X0Y122_I),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000011100000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f000f110f55)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005555e000c000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaabbbbbbbbbbbb)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222000023220000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaabfbfbf)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4044c0004050c0f0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0f070f07)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3020002000003030)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333300505050)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff05ff00ff)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00007777)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000500000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ab00ffffffff)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.I4(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaa888a888a888)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeefe000000f0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.I4(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcdcdcdcdcdcdcc)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_DO6),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f100000000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000220000002000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I1(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddddddddddc)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fffe0000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I5(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050555550505544)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_DO6),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00000000131313)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h080d0000c8dd4000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5d5c5c0ffffc5c0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h11111111ffff1f11)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000044440f020f00)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff33ffff)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffe)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f100000011)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0008000f333a222)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303030355fd00fc)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h73ff73ff50ff50ff)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f300f351510051)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7fffffff3fff3)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2fff2f2fffffff2)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbfffff)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aafffffcfefcfe)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000031113333)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y127_IOB_X0Y127_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fe00aa00ff00aa)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(LIOB33_X0Y121_IOB_X0Y122_I),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabafafa30baf0fa)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f000f888f)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h008a008a0000008a)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000505500001011)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_CO6),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_CO6),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdddf)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I1(CLBLL_L_X2Y116_SLICE_X1Y116_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a00000022000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3ff0000bbff0000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0affceffceffce)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffeefffcfffeff)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I3(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_CO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000101cc00dc00)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002000000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.I1(CLBLL_L_X2Y116_SLICE_X1Y116_BO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3131f5f5ccc00000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000f00040005)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_DO6),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf555f000f7fff0cc)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa00fafafa00fa32)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff880f0a0f08)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccf888f000f000f)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000005050d0dcdcd)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(1'b1),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333000033333030)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(1'b1),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbaaaaaaaa)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_BO6),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa000c040800)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_BO6),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f1f0f5f5f0f0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffcfaa88ffcc)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcdcdcdffffcdcd)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_DO6),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(1'b1),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88ff80f0fffff0f0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffa0f080c0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_DO6),
.I3(RIOB33_X105Y119_IOB_X1Y120_I),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aabb0000afbf)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(RIOB33_X105Y119_IOB_X1Y120_I),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001100100010)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3733ffff3333)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_DO6),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f0c3f3f3f0d)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffeffeefffe)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3f373f3f)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.I1(LIOB33_X0Y121_IOB_X0Y121_I),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf555c444ffffcccc)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I5(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050511111111)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0dfd0dfd00000300)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaaaaae)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(RIOB33_X105Y115_IOB_X1Y115_I),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cf0000000a00)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff8c88cccc)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f3f30f000c00)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heefeeefefefefefe)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeea0e0aaeeaaee)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0cff0cff4cff0c)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000101ffe8ff80)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff8880)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555700000003)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffff00ec00ee)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22ff22ff55550000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaacc8888000000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(1'b1),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00aaf0fff0fa)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(1'b1),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfcfffffdfcfdfc)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b03030b0bb3033)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y124_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc0000cdcc0000)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0545050505050507)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y115_IOB_X1Y115_I),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafafafaf8f)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.I3(RIOB33_X105Y113_IOB_X1Y114_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y115_IOB_X1Y116_I),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3331331131311111)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000ff0affaa)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I1(1'b1),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y124_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y126_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y127_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_BO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X2Y132_SLICE_X0Y132_AO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X2Y127_SLICE_X0Y127_AO5),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_AO6),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X2Y125_SLICE_X0Y125_AO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y127_SLICE_X0Y127_AO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLL_L_X2Y130_SLICE_X0Y130_AO5),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_AMUX = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_AMUX = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_AMUX = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_AMUX = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D = CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_AMUX = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_BMUX = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_DMUX = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_AMUX = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_BMUX = CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_CMUX = CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_AMUX = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_BMUX = CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AMUX = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_AMUX = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_AMUX = CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_BMUX = CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D = CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D = CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B = CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D = CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_AMUX = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A = CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B = CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C = CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D = CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B = CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D = CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A = CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B = CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D = CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D = CLBLL_L_X2Y130_SLICE_X0Y130_DO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_AMUX = CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A = CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B = CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D = CLBLL_L_X2Y130_SLICE_X1Y130_DO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A = CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B = CLBLL_L_X2Y132_SLICE_X0Y132_BO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C = CLBLL_L_X2Y132_SLICE_X0Y132_CO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D = CLBLL_L_X2Y132_SLICE_X0Y132_DO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A = CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B = CLBLL_L_X2Y132_SLICE_X1Y132_BO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C = CLBLL_L_X2Y132_SLICE_X1Y132_CO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D = CLBLL_L_X2Y132_SLICE_X1Y132_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C = CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D = CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A = CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B = CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C = CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D = CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AMUX = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_AMUX = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_BMUX = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AMUX = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_AMUX = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_AMUX = CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AMUX = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_AMUX = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_CMUX = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AMUX = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_AMUX = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_AMUX = CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_AMUX = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_AMUX = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_BMUX = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_AMUX = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_BMUX = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_DMUX = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_AMUX = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_BMUX = CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_AMUX = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_AMUX = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_AMUX = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_BMUX = CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_AMUX = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_AMUX = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_AMUX = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A3 = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A5 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A1 = CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A2 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A3 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A4 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A5 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A4 = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A1 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A1 = CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A2 = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A3 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A4 = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A6 = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A1 = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A2 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A3 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A5 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B6 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A1 = CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A6 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B4 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A3 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A5 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B1 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B4 = 1'b1;
endmodule
