module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AMUX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_AO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_A_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_BO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_BO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_B_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_CO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_CO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_C_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_DO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_DO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X54Y127_D_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_AO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_AO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_A_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_BO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_BO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_B_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_CO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_CO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_C_XOR;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D1;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D2;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D3;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D4;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_DO5;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_DO6;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D_CY;
  wire [0:0] CLBLL_L_X36Y127_SLICE_X55Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CLK;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C5Q;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CLK;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D5Q;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B5Q;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B5Q;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CLK;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CLK;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C5Q;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A5Q;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B5Q;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CLK;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D5Q;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A5Q;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CLK;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A5Q;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5Q;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D5Q;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C5Q;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C5Q;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5Q;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5Q;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A5Q;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AMUX;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BMUX;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DMUX;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AMUX;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C5Q;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CLK;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A5Q;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B5Q;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CLK;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B5Q;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A5Q;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CLK;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CLK;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CLK;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CLK;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AMUX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CE;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_SR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CLK;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CLK;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CLK;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CE;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CLK;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_SR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CLK;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5Q;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D5Q;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D5Q;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B5Q;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CMUX;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CMUX;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5Q;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5Q;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_XOR;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A1;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A2;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A3;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A4;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_AO5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_AO6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A_CY;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_A_XOR;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B1;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B2;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B3;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B4;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_BO5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_BO6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B_CY;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_B_XOR;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C1;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C2;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C3;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C4;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_CO5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_CO6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C_CY;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_C_XOR;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D1;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D2;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D3;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D4;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_DO5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_DO6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D_CY;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X162Y139_D_XOR;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A1;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A2;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A3;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A4;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_AMUX;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_AO5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_AO6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A_CY;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_A_XOR;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B1;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B2;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B3;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B4;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_BO5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_BO6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B_CY;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_B_XOR;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C1;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C2;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C3;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C4;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_CO5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_CO6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C_CY;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_C_XOR;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D1;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D2;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D3;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D4;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_DO5;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_DO6;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D_CY;
  wire [0:0] CLBLM_R_X103Y139_SLICE_X163Y139_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AMUX;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AMUX;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_AO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_AO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_BO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_BO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_CO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_CO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_DO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_DO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_AO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_BO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_BO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_CO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_CO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_DO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_DO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AMUX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AMUX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BMUX;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CMUX;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A5Q;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C5Q;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D5Q;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D5Q;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5Q;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C5Q;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BMUX;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B5Q;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CE;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_SR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A5Q;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CLK;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CLK;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CE;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CLK;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_SR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CLK;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CLK;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_BO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CLK;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_DO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AMUX;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CLK;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_DO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CLK;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_DO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A5Q;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AMUX;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AX;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BMUX;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CLK;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_DO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CLK;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_DO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AMUX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BMUX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CE;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CLK;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CMUX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_SR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BQ;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CLK;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_DO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CLK;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CMUX;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DMUX;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CLK;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BQ;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CLK;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CLK;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CLK;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CMUX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CLK;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CLK;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CLK;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CLK;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CMUX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CLK;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_CO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_DO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_AO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_AO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_BO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_CO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_DO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_DO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_AO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_AO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_BO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_DO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_DO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_AO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_AO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_BO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_DO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_BO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_BO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CLK;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_DO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_DO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_BO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_BO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CLK;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_DO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_DO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_AO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_AO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_BO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_BO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_CLK;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_CO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_CO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_DO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_DO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_AO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_AO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_BO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_BO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_CO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_CO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_DO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_DO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CLK;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AQ;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CLK;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CLK;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CLK;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AQ;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BQ;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CLK;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_DO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_BO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CLK;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_DO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CLK;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CLK;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CLK;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A5Q;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AMUX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DMUX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5Q;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C5Q;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D5Q;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A5Q;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5Q;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5Q;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5Q;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B5Q;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CE;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc330000cccc)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_DO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffdfffffffcf)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffefffcfffff)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfdffffffdd)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I4(CLBLM_R_X3Y130_SLICE_X2Y130_BQ),
.I5(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_CO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_DO5),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_AO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_CO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_DO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaccaacc)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_DLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_CLUT (
.I0(RIOB33_X105Y127_IOB_X1Y127_I),
.I1(CLBLL_L_X4Y123_SLICE_X5Y123_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f06600cc00)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I1(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_DO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88d888d888d888d8)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_D5Q),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_CO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005f5fff33ff33)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_DLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000000fff0fff)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaf0005aaae0004)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_DO5),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I5(CLBLL_L_X4Y124_SLICE_X4Y124_CO6),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaa040033ff33ff)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_BO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_DLUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_A5Q),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa088880000)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_CLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I1(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y127_IOB_X1Y127_I),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5f00a000)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_BLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_DO6),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0048484848)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_ALUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_DO6),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_CO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aafff0f088cc)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_CQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_BLUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_CQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AQ),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000dddc1110)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_DO5),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_BO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05ff0fff55ffffff)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff135f80008000)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_CLUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_A5Q),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14aa00be14aa00)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_CO5),
.I3(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1c0e2c0d1c0e2c0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X4Y126_AO6),
.Q(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.Q(CLBLL_L_X4Y126_SLICE_X4Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f7fffff7f7ffff)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafef000000cc00cc)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_B5Q),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_C5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9fc090cf0f00000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_BLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.I4(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3ffaaaac000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_ALUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_B5Q),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X5Y126_AO6),
.Q(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X5Y126_BO6),
.Q(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdcff50dcdc5050)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_BO5),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300000013000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_B5Q),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccff00f0f0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_B5Q),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccf0ccaacca0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y123_SLICE_X6Y123_DO6),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_BO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_CO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f0aaaa)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3030f0f0ff00)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_CLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_DQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cf000fc0c)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc005acccc005a)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_DO6),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_DO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0ead5aaffaaff)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_DLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_B5Q),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_A5Q),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088f022f022)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_CLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff030003ff030003)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_C5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcdecccc30120000)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_ALUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.I5(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_BO5),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_CO5),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_DO5),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_BO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_CO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_DO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cafa0afa0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_DLUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I2(CLBLL_L_X4Y124_SLICE_X4Y124_B5Q),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500ecececec)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_DO6),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3ffaaaac000)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_ALUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_BO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_AO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030123030303030)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_DLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_B5Q),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_A5Q),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfffbffbbbb0000)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacaca0000aa00)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f000f000)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_DO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h005000ff00500050)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_DLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I1(1'b1),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202000002020f00)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_CLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_BQ),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffefee)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_BLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_DO6),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_CO6),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_AO6),
.I5(CLBLM_R_X3Y129_SLICE_X3Y129_CO6),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005500ff307530)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_CQ),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_DQ),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000aacc)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_DLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_A5Q),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffeffffff)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_BLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeffeffffff)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000003300f3f0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.I2(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444f4f4ff44fff4)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_CLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_DO6),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_BO6),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_CO6),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_AO6),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_BO6),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000222200f022f2)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3030ff30)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_CO6),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffcf)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_CO6),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_DO6),
.I3(CLBLM_R_X5Y129_SLICE_X7Y129_DO6),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_DO6),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_BO6),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fcf0eeaafefa)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_BLUT (
.I0(LIOB33_X0Y65_IOB_X0Y66_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I2(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_AO6),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff2)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_ALUT (
.I0(LIOB33_X0Y65_IOB_X0Y66_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AO6),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_AO6),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_CO6),
.I5(CLBLM_R_X5Y129_SLICE_X7Y129_DO6),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccfceefeeefe)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_DLUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CO6),
.I2(LIOB33_X0Y67_IOB_X0Y68_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff75ffff3030)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.I2(LIOB33_X0Y67_IOB_X0Y67_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffe)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_BLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_DO6),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_BO6),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_CO6),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_CO6),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_CO6),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffe)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_DO6),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_DO6),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_DO6),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f000c0c0f0c)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f35073f0f05050)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f3fbf0fa)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_CO5),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffba)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_DO6),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_BO6),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AO6),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_CO6),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77ff33ff55ff00)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_DLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_DO6),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_DO6),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_CO6),
.I4(CLBLL_L_X4Y132_SLICE_X4Y132_DO6),
.I5(CLBLL_L_X4Y132_SLICE_X4Y132_BO6),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffa0ec)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_CO6),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_CO6),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff3fbf0fa)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_ALUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_DO6),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_DO6),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222222222222)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_DLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff30ffffff30ff30)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_CO6),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f550f00dfddcfcc)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_BLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_BO6),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_AO6),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000200000)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000ffe5)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7777ffff77f7)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_CLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7ffffffffbffff)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5eff7fffffff7f)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaffbababaffbaba)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_DLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_CO6),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd0000ddfd00f0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(LIOB33_X0Y71_IOB_X0Y71_I),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_C5Q),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00c00008)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_CO6),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfdffffff)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7fffffff5f)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_DLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_CO6),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.I5(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808000000080000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_BLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffffff00ffff)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfcffff3074ff)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffff0000cc00)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y127_SLICE_X54Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y127_SLICE_X54Y127_DO5),
.O6(CLBLL_L_X36Y127_SLICE_X54Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y127_SLICE_X54Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y127_SLICE_X54Y127_CO5),
.O6(CLBLL_L_X36Y127_SLICE_X54Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y127_SLICE_X54Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y127_SLICE_X54Y127_BO5),
.O6(CLBLL_L_X36Y127_SLICE_X54Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055000000550000)
  ) CLBLL_L_X36Y127_SLICE_X54Y127_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_BQ),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y127_SLICE_X54Y127_AO5),
.O6(CLBLL_L_X36Y127_SLICE_X54Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y127_SLICE_X55Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y127_SLICE_X55Y127_DO5),
.O6(CLBLL_L_X36Y127_SLICE_X55Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y127_SLICE_X55Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y127_SLICE_X55Y127_CO5),
.O6(CLBLL_L_X36Y127_SLICE_X55Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y127_SLICE_X55Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y127_SLICE_X55Y127_BO5),
.O6(CLBLL_L_X36Y127_SLICE_X55Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y127_SLICE_X55Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y127_SLICE_X55Y127_AO5),
.O6(CLBLL_L_X36Y127_SLICE_X55Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50aa00eeeeffff)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_A5Q),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffee00ee)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ee44)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccaaccf0cca0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_CO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003321212121)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_DLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_D5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3f3d1d1)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ff33cc00)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000eeec2220)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_CO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_DO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbba1110bbba1110)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f2f1f201020102)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cccc0ff0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0cfcfc0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_CO6),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_DO5),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_CO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ffcc00cc)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeeee00004444)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f08888)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000eee0eee0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_BO6),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0e)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_DLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_A5Q),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.I2(CLBLM_L_X12Y128_SLICE_X17Y128_BQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_DO6),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_D5Q),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafe)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc8ccccccc40cc00)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_BLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_D5Q),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacac0f0f0fff)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1441822814418228)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_CQ),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333300033332200)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_CLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_CO6),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002fffdfcfffcff)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefceefceefceecc)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_DO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff500050ff500050)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e0e0e0e0e0e0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_CLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fe0ef000f000)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_D5Q),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_CO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffeaff50ff40)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_DQ),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_CO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000affa0550)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_CO6),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_A5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff660066)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_BLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff03ff0c0003000c)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_BO6),
.I5(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_DO5),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0aa3a3a0a0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_DLUT (
.I0(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_C5Q),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f40104f1f40104)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habae0104aeae0404)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00af05fa50)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_R_X13Y125_SLICE_X19Y125_BQ),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_BO6),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_AO5),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00d00000f000f)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000a0aa0a0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_DO6),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_DQ),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcc0300cfcc0300)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0f0ccf0cc)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_ALUT (
.I0(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000efff00000fff)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_DLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_CO5),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f000ee00ee00)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cff5f00500)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_BLUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_B5Q),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaeeea55504440)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_BO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669966)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0f0808080f0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_CO6),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1b1a0a0b1b1a0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88dd88ddd8d8)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X11Y123_BO6),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_DLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcc0a0000f0f0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000050055005)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffeaaa51554000)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I5(CLBLM_L_X12Y128_SLICE_X17Y128_BQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_DO6),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I4(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_BO6),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0c0a080000aaaa)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ea40aa00ea40)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_CQ),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000abaa0100)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_CO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_DO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfc00fc)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_DLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_DQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffbe55445514)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fc0cfc0c)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3330fff0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_ALUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_CO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_DO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heecceecc22002200)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_C5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffac00acffac00ac)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefaee50445044)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff33cc00fc30)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_BO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_CO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_DO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd8ffd800d800d8)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_DLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0aaf0ccf0aa)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_CLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f4f405050404)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y130_SLICE_X15Y130_CQ),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_DQ),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88d8ddddd8d8)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000c000808)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_DLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_DO6),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffefffffff)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_DQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdd00aa00aa)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_BLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff320032ff320032)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_C5Q),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I2(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_CO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_DO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044aaea0040)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0aca0ac)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fefe00000e0e)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100ddcc1100)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_DQ),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_CO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fe32fe32)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_D5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_DQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54ae04fe54ae04)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf8fdf80d080d08)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_DQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff505050505050)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000000)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefedcdc32321010)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_CO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505000505000000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_DLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I1(1'b1),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_DQ),
.I5(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaaa00550000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I5(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f60606f0f00000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00d2d2ff000000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_ALUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_BO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0000b3a0b3a0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_A5Q),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04ae04ae04ae04)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3030aaaa3030)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaacccc)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_C5Q),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0f0aa0000f0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_B5Q),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000030303030)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_D5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000a800a8)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f044f044)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccfacc50)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff540054ff540054)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff5000550050)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_CO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_DO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f033003300)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c0c0cccc)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0dd88f0f05500)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I3(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0ccaaaa00cc)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa0088ffaaffbb)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_DLUT (
.I0(CLBLM_R_X13Y121_SLICE_X18Y121_BO6),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_D5Q),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7272723327272733)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_D5Q),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ee22ff33)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff32ff3200320032)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_ALUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00ee00ff00ff)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_DLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_A5Q),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdc001033303330)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ff000000)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_DLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f99959995)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_CLUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f80808cfc0cfc0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I4(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaafcaa00)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_B5Q),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_DQ),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd888dd8dd88dd88)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.I4(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cc993369c369c3)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_BQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_CQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22020000aaaa8888)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa30aa33aa30)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7fffffff7ffff)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccfccc0c)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fc30fc30)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31ec20dd11cc00)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc048800cc008800)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_DLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f000ee00ee00)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_CLUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff00decc5a00)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaf0f0cc00)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_ALUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_A5Q),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_DLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000033003300)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aa30aa30)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00fafa)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_ALUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00aaaaaaa8a8)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_DO6),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa800a8a8a8a8a8)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000eee0eee0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000c800c8)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_DLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_CO6),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_A5Q),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_DO6),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef00e00ee00ee00)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_DQ),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf2faf20a020a02)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050005)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_DLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdf111100000000)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa88aa88fafa5050)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf011f022f011f022)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_ALUT (
.I0(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafa)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_DLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_C5Q),
.I3(1'b1),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffc)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000003535353a)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_BLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_BO6),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaababa00001010)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_D5Q),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heecfeecceecfeecc)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_DLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfaf80f0c0a08)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_CLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_CO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1c0c0ffcc3300)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_C5Q),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f5f000050500)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.I5(CLBLM_L_X10Y128_SLICE_X12Y128_C5Q),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_DO5),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_DO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2eeee2222)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_DLUT (
.I0(RIOB33_X105Y125_IOB_X1Y126_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff55af05)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I5(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaa00fcfc0000)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_BLUT (
.I0(CLBLM_R_X3Y128_SLICE_X2Y128_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fcfca8a8)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_DO6),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_CO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_DO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5a0f5a0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100f3f3c0c0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_CQ),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefef00e0e0e00)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_BLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_DO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa50fa50)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(1'b1),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_BO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fff00000eeee)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_A5Q),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcf80c08)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.I5(CLBLM_L_X8Y126_SLICE_X11Y126_CO6),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cf000fc0cf000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_CO5),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_BO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5f500ff0033)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ee44d8d8d8d8)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_CQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I3(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafc0a0a0a0c)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_BLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_DQ),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333ff003030)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_BO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005050000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I1(1'b1),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(1'b1),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888b88b8bb8)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_BQ),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fff0ffb0b)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y125_SLICE_X17Y125_B5Q),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfce0302cccc0000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_DO6),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_CO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_DO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0044444444)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55005500)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_A5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef40e04fef40e04)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aa00aaf0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I5(CLBLM_R_X11Y130_SLICE_X15Y130_BQ),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_BO6),
.Q(CLBLM_L_X10Y130_SLICE_X13Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X13Y130_BO6),
.Q(CLBLM_L_X10Y130_SLICE_X13Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.Q(CLBLM_L_X10Y130_SLICE_X13Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X13Y130_DO6),
.Q(CLBLM_L_X10Y130_SLICE_X13Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fe54fa50fa50)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_BQ),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_DO6),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888d8d8d8d8)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_CO6),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0acafafa0aca0a0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_DQ),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202ff0ff202f000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_CO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0000fafa)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0e2e2c0c0e2f3)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_A5Q),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5f40f0f0504)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff44e4000044e4)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hecec2020eeec2220)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_DQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_DQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05aa00ef45ea40)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fdf0f8050d0008)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbffff0f0b0f0f)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_DQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044444444)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e0f00001100)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fdf0f8050d0008)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff5accccff5a)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_CO6),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffccfffe0000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_DQ),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffaa00aa)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(RIOB33_X105Y143_IOB_X1Y144_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0c0c030c)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_CQ),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcffcc10103300)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_C5Q),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500040000)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005454ff001010)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_BO5),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055541154)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_BO5),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00b0f000f0f00000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_DO6),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeaeafffff000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff752000007520)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_ALUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_DQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0fff3f3f3f3)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff01dd10ff02ee2)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_DLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_B5Q),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_AO6),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e40f4ef0b10f1b)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_AO6),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_A5Q),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c000aaaaaaa6)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_BLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_CO6),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa9aaa0000ff00)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_BO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_CO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_DO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888ddd888888888)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_DQ),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00008f808f80)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf8aa88f8fa88aa)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaa603030303)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffff55aaffffaa)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_DLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I4(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fffff0ff0fffff0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I4(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeffffbebeffffbe)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaffaa00aaf0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_ALUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_CO6),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X17Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_DLUT (
.I0(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcffcffffcffc)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff2fff1fff)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_BLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_BO6),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.I5(CLBLM_L_X12Y122_SLICE_X17Y122_CO6),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005454ff005454)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_AO5),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ffff33ccffffcc)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333ccccffcc)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_CQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffcfffef0010)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_BLUT (
.I0(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fafa0a0a)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_ALUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_A5Q),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_BO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0131023201310131)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_DLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_BO6),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fa50aa00ff55)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X17Y123_DO6),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00d5d5ff008080)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0d2f0f0ffffccff)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_ALUT (
.I0(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_AO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_BO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_CO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_DO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccfcfcecec)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_DLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_CO6),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_DQ),
.I3(CLBLM_L_X12Y124_SLICE_X16Y124_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff554400005544)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_CQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_A5Q),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000fcfc)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I3(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00d5d5ff008080)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_AO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_BO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_CO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0407040704070704)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_DLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_A5Q),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I4(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaee00550044)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf00c00fafa0a0a)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_BLUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_AQ),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fe32cc00dc10)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_L_X12Y121_SLICE_X17Y121_DQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_CO5),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_DLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_BO5),
.I3(CLBLM_R_X13Y125_SLICE_X19Y125_BQ),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_CLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_A5Q),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0f0f0f00)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_BQ),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.I3(CLBLM_R_X13Y125_SLICE_X19Y125_BQ),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33333030)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y125_SLICE_X18Y125_AO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_CO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_AO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_BO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y125_SLICE_X17Y125_DO6),
.Q(CLBLM_L_X12Y125_SLICE_X17Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cc00ce02cc00)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_DLUT (
.I0(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_L_X12Y125_SLICE_X17Y125_DQ),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8888800300030)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_CLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I4(CLBLM_L_X12Y125_SLICE_X17Y125_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0010104040)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dc10cc00cc00)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X17Y125_DQ),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_BO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_CO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0110233201012323)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_CQ),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_B5Q),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0aca000ff33ff)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_CLUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I1(CLBLM_R_X13Y126_SLICE_X19Y126_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0c0c0f3c0c0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfddd3111eccc2000)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044aaff0055)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_DO6),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5e4f5e4)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I2(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f2f0f800020008)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaf0aac0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_D5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_BO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_CO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_DO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aaccaac0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_DLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa0faaf0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_CLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ea40f0f0c0c0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_BQ),
.I4(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00fa00fa)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.I1(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X17Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.Q(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X17Y127_CO6),
.Q(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ee00ee00ff00f0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_DLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafcfafcfafcfaf0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_CLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_C5Q),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_CQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0e40000f0e4)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_BLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000b8b8b8b8)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_AO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_BO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_CO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_DO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaf0aac0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_DO6),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888b8bb8b8)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_CLUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffffaaaa)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y131_SLICE_X17Y131_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc0f0cf3f00300)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y130_SLICE_X17Y130_BO6),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_AQ),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_CO6),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X17Y128_AO6),
.Q(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X17Y128_BO6),
.Q(CLBLM_L_X12Y128_SLICE_X17Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000c0c0c0c)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y128_SLICE_X17Y128_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ff00fcfc)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X16Y129_AO6),
.Q(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.Q(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffff)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333303033223322)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I3(CLBLM_L_X12Y124_SLICE_X16Y124_DQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fef0f0000e0000)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_BLUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_DO6),
.I1(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ccccaaaa)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_ALUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.I1(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X17Y129_AO6),
.Q(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.Q(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.Q(CLBLM_L_X12Y129_SLICE_X17Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X17Y129_DO6),
.Q(CLBLM_L_X12Y129_SLICE_X17Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00ba10aa00)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_DQ),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_CQ),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfaaafa11500050)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_CQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0e4f5f5a0a0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I4(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I5(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0aca0aca0aca0ac)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_DQ),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_AO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_BO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_CO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_DO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcccd03030001)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_DLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I4(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0a000affca00ca)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_CLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_CQ),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cac0cacfcac0ca)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_BLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccf0cc00cc5a)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_ALUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_CO6),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.Q(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.R(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7333dd9973cc77cc)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.I3(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5d5f0c0f5f5f0f0)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_BLUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I1(CLBLM_L_X12Y130_SLICE_X17Y130_CO6),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_CO6),
.I4(CLBLM_L_X12Y130_SLICE_X17Y130_AO6),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_CQ),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044004407070707)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_CO6),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_DO6),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc32cc00cc00)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_DLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I1(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_BQ),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafeeaaee05440044)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_CQ),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hececececfff0ff00)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_BLUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_DQ),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_BO6),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaafcaa00aa30)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_CQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y131_SLICE_X17Y131_AO6),
.Q(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0045004500550050)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y131_SLICE_X17Y131_BO5),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f0533333332)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000200)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_BLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I3(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff33aaaaff30)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_DQ),
.I1(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_CQ),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa59aa55aa95)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_DLUT (
.I0(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I5(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333312333333333)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000004)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_AQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0032321010)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_ALUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_A5Q),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_AO6),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_BO6),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_CO6),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4003100f5f5f5f5)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_CQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_DQ),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_DO6),
.I5(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0dfd0dfc0cfc0c)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y132_SLICE_X17Y132_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff030f00ff000f)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_AO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_BO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_CO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c9c3c9c3c9c3c3)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_DLUT (
.I0(CLBLM_L_X10Y130_SLICE_X13Y130_BQ),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.I5(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000bbbbb0b0bbbb)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_CLUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.I5(CLBLM_R_X11Y133_SLICE_X15Y133_CO6),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd755d7550000d755)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_BLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_CO6),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h45cf00cf45cf00cf)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_ALUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.Q(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.R(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y137_SLICE_X16Y137_AO6),
.Q(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0c0dddddddd)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc80cccccc8080)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_B5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_DO6),
.I5(LIOB33_X0Y51_IOB_X0Y51_I),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffcfffffffaf)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X3Y124_AO6),
.Q(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000050005000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.Q(CLBLM_R_X3Y125_SLICE_X3Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11bb11ba10ba10)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_DO6),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_ALUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_BQ),
.I5(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_BO6),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a5a5ff000000)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff9c009cff000000)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaafeaafc00fc00)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_BLUT (
.I0(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_BQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_DQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeccfeccfa00fa00)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_DQ),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X3Y127_DO5),
.Q(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.Q(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.Q(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X3Y127_CO6),
.Q(CLBLM_R_X3Y127_SLICE_X3Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000a8a0a0a0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_DLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_BQ),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088f000f0aa)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_CLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_CQ),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_DO6),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00a8000000a8)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_BLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_CQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00b0b0b0b0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_B5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.Q(CLBLM_R_X3Y128_SLICE_X2Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y128_SLICE_X2Y128_BO6),
.Q(CLBLM_R_X3Y128_SLICE_X2Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_DO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_CO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01144f0f00000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_BLUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I1(CLBLM_R_X3Y128_SLICE_X2Y128_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_B5Q),
.I3(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_BO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfeaffaa15405500)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y128_SLICE_X2Y128_BQ),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I4(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_AO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.Q(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_DO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_CO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_BO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fe540000fe54)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I2(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.I3(CLBLM_R_X3Y128_SLICE_X2Y128_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_AO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.Q(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X2Y129_BO6),
.Q(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_CLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff6000000060)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_BLUT (
.I0(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaeea00000440)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I3(CLBLM_R_X3Y130_SLICE_X2Y130_DO5),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_AO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_BO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h002f0022002f0022)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_DLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020000000000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_CLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00d8d8d8d8)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_BLUT (
.I0(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafffcaaaa0030)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X2Y130_CO6),
.Q(CLBLM_R_X3Y130_SLICE_X2Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X2Y130_AO6),
.Q(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.Q(CLBLM_R_X3Y130_SLICE_X2Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_DLUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0c0c00000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_BQ),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.I4(CLBLM_R_X3Y130_SLICE_X2Y130_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f00100f2f00200)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_BLUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_DO6),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_A5Q),
.I5(CLBLM_R_X3Y130_SLICE_X2Y130_BQ),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3cfaf0aa00aa00)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y128_SLICE_X2Y128_BQ),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I4(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000312000000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I2(LIOB33_X0Y57_IOB_X0Y57_I),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_BQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffffffffaf)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeffffeffffff)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_CO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_AO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_BO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haf00bf33af00af00)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I5(LIOB33_X0Y67_IOB_X0Y67_I),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0c011110000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa03000c00)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X2Y131_SLICE_X1Y131_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3caa00faf0aa00)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_AO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5f5f5f5)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000220000001010)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heffffffffeffffff)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00003c00)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_ALUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I1(CLBLL_L_X2Y131_SLICE_X1Y131_AO6),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f500f0ddfdccfc)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_DLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_AO6),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I2(LIOB33_X0Y59_IOB_X0Y59_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_BO6),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020002000220000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.I2(LIOB33_X0Y59_IOB_X0Y59_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffffffff3fffff)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_BLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbffeffffff)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_ALUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffffffff)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888f888888888)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_CLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff4)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_ALUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_DQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.I3(CLBLM_R_X3Y132_SLICE_X3Y132_BO6),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_CO6),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_CO6),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffff03002000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffffefffff)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0041410000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc8c8c8c8c8c8)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_ALUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_BO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_CO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0a3a0a3)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa03aa0caa03aa0c)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_CLUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_D5Q),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y123_SLICE_X6Y123_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f055f000f0aa)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_BLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaf0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_DO6),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_DO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_BO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_CO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdffd1331f000f000)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_A5Q),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff6600000066)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_BO6),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeaaaaffcc0000)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I5(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffa00fa00fa00)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_BO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_CO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0ffa0a0ecffecec)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I2(CLBLM_R_X3Y128_SLICE_X2Y128_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I5(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0ccaaaaf0f0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_CLUT (
.I0(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f8f8aa00ff55)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_BQ),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_DO6),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88d8ddddd8d8)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff33)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_CO6),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_A5Q),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcff)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_D5Q),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_B5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_A5Q),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_CO6),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fedc3210)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_DLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa20aaaadfdfdfdf)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_DQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3c0b8b8b8b8)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdecc1200fccc3000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_C5Q),
.I1(CLBLM_R_X3Y130_SLICE_X2Y130_A5Q),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_C5Q),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_C5Q),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_C5Q),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_C5Q),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_D5Q),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_DO6),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_C5Q),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_A5Q),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffee)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_ALUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_A5Q),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_B5Q),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_CO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5010ffffffff)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e0e0ff00eeee)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0fc00fc00)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044eeee4444)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080808000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_A5Q),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff3369969669)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf088f0fff0cc)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaa0ccccfff0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_DO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fa50ee44ee44)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_A5Q),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acacaca0a0a0a0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_A5Q),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e4e4ff00e4e4)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdc5050dcdc5050)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaaaaaaa)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_C5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_D5Q),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5555cccc0000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_DQ),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf8fdf80d080d08)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0f0ff00)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_CQ),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_CO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaafaaabffffffff)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_B5Q),
.I3(LIOB33_X0Y53_IOB_X0Y53_I),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_A5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff800000008000)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_CLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_A5Q),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0cc00cc00cc00)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_A5Q),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_C5Q),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_B5Q),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefcc2300efff2333)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_ALUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I5(LIOB33_X0Y53_IOB_X0Y53_I),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_CO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000b000b00080008)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_DLUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0cfcfc0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccffaaaacc00)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeba5410feba5410)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0aafa00f0aafa)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_C5Q),
.I3(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f33330f0f0000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_BO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f500f0ddfdccfc)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_BLUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_AO6),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffcfffdfdfcfc)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_CO6),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AO6),
.I3(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h03030b0b00000a0a)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff22ffffff2222)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_AO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_DO6),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c69963cc39669)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaaafafffafa)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I1(1'b1),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0affceff0a0acece)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_B5Q),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_DO6),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_CO6),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_BO6),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_BO6),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I5(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0f00cfcc)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_DQ),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_BO6),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00004f4400004f44)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h005500000c5d0c0c)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdfcfcf00550000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefffefffefefefe)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_DO6),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_CO6),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_CO6),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_DO6),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_BO6),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffffffffff)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080008000a00000)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BO6),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabababaffffbaba)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_DLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb00bb00bb00fbf0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb8ffb800b800b8)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_A5Q),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f1f01100)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_A5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DO6),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_BO6),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_DO6),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_AO6),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_DO6),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_CO6),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_BO6),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_AO6),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_AO6),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffffffaaaaffff)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff3bff0a)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_CO6),
.I4(LIOB33_X0Y65_IOB_X0Y65_I),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_BO6),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffffffefe)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_CLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_CO6),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_DO6),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_DO6),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000000)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_BLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_CQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033507300005050)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_ALUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000003120)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffae)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_BLUT (
.I0(CLBLM_R_X5Y133_SLICE_X6Y133_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_DO6),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_CO6),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_ALUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_CO6),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_AO6),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeff00004400)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_BLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h40400000fcffffff)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_ALUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400040)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaaabfffbfbf)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_CLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_AO6),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbfffffff)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_DO6),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_CO6),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f8f0fa)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5ffffffaffffff)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(1'b1),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaaee00440044)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454feaa5400)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_C5Q),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff33ff33)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffffffffffff)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11ba10bb11ba10)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf5fffff8f0ffff)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I3(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaafe00cc00fc)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_CQ),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaaaaaba10000010)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I5(CLBLM_L_X12Y124_SLICE_X16Y124_DQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000eefdaaf5)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb33333333)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff080800000808)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c5c5c0c0caca)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_B5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffe000e0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff78f0000078f0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff01a801ff00aa00)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0aaf0ccf088)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_CO6),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff00fcfc0000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffaa)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_DLUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y125_SLICE_X17Y125_B5Q),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5fffffffffff)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_CLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I4(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I5(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000e000e0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_DQ),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33303330)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc8ccc0c0d1c0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ccccecff)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.I2(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_CO6),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h05050505afafafaf)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccf0cca0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aaccaacc)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_A5Q),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c000cccaaccaa)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_CLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0012121212)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff00fafa0000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_CO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033393333)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_A5Q),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I5(CLBLM_R_X3Y125_SLICE_X3Y125_AQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ce020a0a0a0a)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_CLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaff0f0f)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DQ),
.I1(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I2(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007474ff00f0f0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3bffbbff0a0aaaaa)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffffffffff)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a00000055ff55ff)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa3cf0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeae0030eeee0000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaf00afff8c008c)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f00000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00faccccfafa)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_B5Q),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100010)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_DLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_CO6),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_DO6),
.I3(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_CO6),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacafa0acacafa0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_CLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_C5Q),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf707ff0fff0fff0f)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_BLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_B5Q),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_C5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000440000)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_ALUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_B5Q),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_CO6),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h13135f5f0000ff00)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_CLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa3c3c)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_CO5),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4a0b1f5a0a0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_BO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_CO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d888d88c0c00000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_B5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0af3f00300)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0b1f5e4a0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_C5Q),
.I3(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88ddd8ddd8)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_DO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf800fa00fc00ff00)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_DO6),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_DO6),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffffff)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_CLUT (
.I0(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c5cac5ca)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_BLUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00f0ccccaafa)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_DO6),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_BO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_CO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_DO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffaaaa00f0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cafafa0a0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_CLUT (
.I0(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaaee00440044)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcdddc11101110)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_CO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hba10ba10fe54ba10)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf5fc000c050c)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccffcc00)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0ccf0cc)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0affffff0aff0a)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_DO6),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111111111101110)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e4e4ff00e4e4)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ba10c0c0c0c0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f0000000c000c)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_DQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f3bbfb00f0aafa)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_BO6),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77335500f7f3f5f0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haabb0011aaee0044)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_DO6),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaf0aaf0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef0fef0ee00ee00)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_CQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccee0000)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_BLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888dd88d8d8d8d8)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000312000003120)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfafffffbbaa)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_CLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_BO6),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_CO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303010f0f0f050)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_BLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554111055541110)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00ccaaeeaaee)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004400000050)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfffeffff)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff55e4e4e4e4)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeffffaaeeaaee)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_AO6),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_DQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.I5(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaeefafe)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0aa33aaf0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.I5(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeefffe)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_AO6),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_AO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_CO6),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_BO6),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000e04)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000cc505050dc)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000044444444)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_B5Q),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222ff22ff22)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.I2(1'b1),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfafa0c0c0a0a)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_A5Q),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I5(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y130_SLICE_X2Y130_A5Q),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000fc0cf000)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_DQ),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_C5Q),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000fcfcf0f0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffbb)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(1'b1),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaf0aaccaaf0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_ALUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I1(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_AO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h555f5fff555f5fff)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_CLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcbcbebeb30305252)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_B5Q),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcbcbefef41418181)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_B5Q),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h02000000eccccccc)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_DLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fff5000000f5)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000008822)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccfacc00cc00)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0e2e2f3f3)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_CO6),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00ff50af00)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1013131010101313)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_D5Q),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.I4(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000447700007447)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_AO6),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I4(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f708ffff3333)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_DO6),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I5(CLBLM_R_X11Y123_SLICE_X15Y123_BO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050045405550151)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_CLUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_AO5),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_BO5),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc9c0fff0fff)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaff00bf40)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_BO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_CO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0131013101310131)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000f5f5)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff33f0f0aa22)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ffcc3300)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_D5Q),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669966)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_DLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969669699696)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_CLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a5005a005a00a5)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_BLUT (
.I0(CLBLM_R_X11Y122_SLICE_X15Y122_DO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_CO6),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_BO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffff55aaffffaa)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_D5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_BQ),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_B5Q),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000055445544)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc50cc55cc50)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6fffff6f6fffff6)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_D5Q),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200002211000011)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_CLUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0202fefd0101fd)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_BLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_BO5),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0021000000840000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_A5Q),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BO6),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_DO6),
.I4(CLBLM_R_X11Y123_SLICE_X15Y123_CO6),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_CO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0b0f00000c000)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_DLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_DO6),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330033ff000000)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_B5Q),
.I5(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ff0033)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc50cc55cc50)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000044)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d11111d1d11d1d)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_BLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88d888dd88d8)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_CO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffcc)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_BQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_DQ),
.I5(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaccaacc)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cac0ff00aa00)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_BLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I1(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdd0011ccee0022)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_ALUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.I5(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_BO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_CO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h99999a9a99999a9a)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_BQ),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0af808ff0ffc0c)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y124_SLICE_X16Y124_CQ),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44aa00aa00)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000001680168)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_ALUT (
.I0(CLBLM_R_X11Y125_SLICE_X15Y125_DO6),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_BQ),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_D5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_CO5),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_DO5),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_CO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_DO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaa00aaaaf0f0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_DLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_C5Q),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f00500f404f404)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0c0f0c0f0c0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_CQ),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_A5Q),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00a8a8)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_BO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_DO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000010001000)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88bb88888888)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_A5Q),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afaca0a0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_BLUT (
.I0(CLBLM_R_X13Y126_SLICE_X19Y126_CQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0cfc0c0cfc0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_DO5),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_DO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05aa00dd88dddd)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_DQ),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_BQ),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0f5a0f5a0a0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.I5(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ee00ee00ee00)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_DQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccaaccaaf0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_ALUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_DO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00cc00c0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_DLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ee44aa00ff55)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_DO6),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc4ffc400c400c4)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_D5Q),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcdddc11101110)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_BO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_BO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000a800a8)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_DLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0f0f0000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_CLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_CO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0f0cc)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_BLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfaccfaccfacc00)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_D5Q),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_DQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_DO5),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_BO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002222dc10dc10)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_DQ),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_CQ),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfc0030e2e2e2e2)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccffcc00ccaa)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I1(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_BQ),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbb8b8b8b8)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_CO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff0f)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_CQ),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I5(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa003300cc)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_CLUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y129_SLICE_X14Y129_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cca0f0f0a0a0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_BLUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_DQ),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_B5Q),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccfff0ff00)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X15Y129_BO6),
.Q(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_CQ),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I5(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_CLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_BQ),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_DO6),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_DO6),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_DO6),
.I5(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff4400550044)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffb00fbffff00ff)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_A5Q),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_BO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_CO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00ffe0ffe0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_R_X11Y130_SLICE_X14Y130_DQ),
.I3(CLBLM_L_X8Y123_SLICE_X11Y123_CO6),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f033003300)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_DQ),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccf0f0ff00)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_BLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f044f044)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X15Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X15Y130_BO6),
.Q(CLBLM_R_X11Y130_SLICE_X15Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X15Y130_CO6),
.Q(CLBLM_R_X11Y130_SLICE_X15Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f044221144)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_CQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_CQ),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_CQ),
.I4(CLBLM_R_X11Y130_SLICE_X15Y130_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f000f000f303)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_CO5),
.I5(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfceeee00302222)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_ALUT (
.I0(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I4(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I5(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.R(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_A5Q),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.R(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdd1d1d3322e2e2)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_DQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333373733373)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefefe00f00000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.Q(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a999a9999999999)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808101008881000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa000000005500)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fbfb0b0b)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_DO5),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_BO6),
.Q(CLBLM_R_X11Y132_SLICE_X14Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X14Y132_AO6),
.Q(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00fa50fa5)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_DLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0037ffff0037ffff)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_DQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h48cc48cc0c000c04)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_DO6),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7030773370307733)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_ALUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_DO6),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_CQ),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X15Y132_AO6),
.Q(CLBLM_R_X11Y132_SLICE_X15Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.Q(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cdefffff)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_DLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c000c000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_CLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9909ff0f0000ff0f)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_DO6),
.I1(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h45cf45cf00cf00cf)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.I4(1'b1),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.R(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777777777577)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333200f000f5)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_BLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf0045ff755530af)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_B5Q),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_B5Q),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3133313330333333)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_DLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccec33033313)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_CLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000a0a)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_BLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_CQ),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c022332233)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_BO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4b4a5a5b4a5a5a5)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_CLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_CO6),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I5(CLBLM_R_X11Y133_SLICE_X15Y133_BO6),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000fccff0c0f)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_A5Q),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_CO6),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffb0000fffb)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y132_SLICE_X14Y132_A5Q),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5044004400440044)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_BO6),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_CQ),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(RIOB33_X105Y127_IOB_X1Y128_I),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.Q(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fffcfc0c0c)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y121_SLICE_X18Y121_AO6),
.Q(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff000f000f)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_DO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hececececececfcfc)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_CQ),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_CO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff4040bfbf)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y124_SLICE_X17Y124_CQ),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_BO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcf0f0ccdc0050)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_DQ),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_CO6),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_AO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y121_SLICE_X19Y121_AO6),
.Q(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_DO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_CO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_BO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdec3120ddcc1100)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I4(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_AO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X18Y122_AO6),
.Q(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X18Y122_BO6),
.Q(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I3(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_DO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33333303)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_DO6),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_AO5),
.I4(CLBLM_R_X13Y122_SLICE_X18Y122_DO6),
.I5(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_CO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaafafa44005050)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_BO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0fffffeeee)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_ALUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I1(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_AO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X19Y122_AO6),
.Q(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X19Y122_BO6),
.Q(CLBLM_R_X13Y122_SLICE_X19Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaca3a0afaca3a0a)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_CQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I3(CLBLM_R_X13Y122_SLICE_X19Y122_CO6),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_DO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333323333)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_CLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I2(CLBLM_R_X13Y122_SLICE_X18Y122_DO6),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_DO6),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_BQ),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_CO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffee00cc00ee)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_BLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_R_X13Y122_SLICE_X19Y122_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_A5Q),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_BO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cc55cc00cc55)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_ALUT (
.I0(CLBLM_R_X13Y122_SLICE_X19Y122_DO6),
.I1(CLBLM_R_X13Y122_SLICE_X19Y122_BQ),
.I2(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_AO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_BO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_CO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_DLUT (
.I0(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5e4a0a0f5e4)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_CQ),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555f0f04444)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_BQ),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffe4440000e444)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_CQ),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_BO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd888d888d888d8)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.I2(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I4(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaffeaaa40554000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I4(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y124_SLICE_X18Y124_BO6),
.Q(CLBLM_R_X13Y124_SLICE_X18Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y124_SLICE_X18Y124_AO6),
.Q(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y124_SLICE_X18Y124_CO6),
.Q(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff8080ffffffff)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_DLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_DO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0e4a0b1a0)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_CQ),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_DO6),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_BQ),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_CO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc5000000f0f)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_BO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_CQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_A5Q),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_AO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y124_SLICE_X19Y124_AO6),
.Q(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_DO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_CO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_BO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0ffaa00c000aa)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_ALUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_BQ),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_AO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.Q(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.R(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002a0000002aaa)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_CLUT (
.I0(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h10000000a0000000)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_BLUT (
.I0(CLBLM_L_X12Y125_SLICE_X17Y125_AQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_BQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_BQ),
.I4(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5fa00aa00aa)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_ALUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_A5Q),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I3(CLBLM_L_X12Y125_SLICE_X17Y125_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_AO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y125_SLICE_X19Y125_AO6),
.Q(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y125_SLICE_X19Y125_BO6),
.Q(CLBLM_R_X13Y125_SLICE_X19Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_DO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_CO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y125_SLICE_X19Y125_BQ),
.I2(CLBLM_R_X13Y124_SLICE_X18Y124_A5Q),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_BO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeec0cceaaec00c)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_CO5),
.I2(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I4(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_AO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.Q(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_BO6),
.Q(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000050000000100)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_DLUT (
.I0(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I1(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I4(CLBLM_L_X12Y125_SLICE_X17Y125_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb888805000500)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_CLUT (
.I0(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_A5Q),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0b1a0e4e4)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_DQ),
.I3(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_CO5),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff00ffe0ffe0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.I4(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X19Y126_AO6),
.Q(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X19Y126_BO6),
.Q(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y126_SLICE_X19Y126_CO6),
.Q(CLBLM_R_X13Y126_SLICE_X19Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffc800c8)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_CLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_R_X13Y126_SLICE_X19Y126_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ff33ff33ee22)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_BLUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I5(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff010001ff100010)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.I2(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_AO5),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.Q(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.Q(CLBLM_R_X13Y127_SLICE_X18Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003300000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555575757575)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b888b888b888b88)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfecccc30320000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_BLUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_ALUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_AO6),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_BO6),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_DO6),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faafcaa00aa00)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_DLUT (
.I0(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f011f055f044)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_CQ),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I5(CLBLM_R_X13Y129_SLICE_X19Y129_BO6),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0a0a0a0a)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_BLUT (
.I0(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffba5510ffbe5514)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_BO6),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.Q(CLBLM_R_X13Y128_SLICE_X19Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y128_SLICE_X19Y128_BO6),
.Q(CLBLM_R_X13Y128_SLICE_X19Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h202020a000000000)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_DLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5511440055114400)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_CLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_AQ),
.I2(1'b1),
.I3(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I4(CLBLM_R_X15Y129_SLICE_X20Y129_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0c00000f0c)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y129_SLICE_X19Y129_AO6),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.I3(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3f2f20f030202)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I1(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020a0a005040000)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_DLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haffaaffaafbeaffa)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_CLUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I4(CLBLM_R_X13Y129_SLICE_X18Y129_DO6),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff50d8000050d8)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_BLUT (
.I0(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff440044ffe400e4)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_ALUT (
.I0(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_CQ),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fdf0fdfff2fff2)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I1(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5aaa55aa59aa55)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_CLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_AQ),
.I1(CLBLM_R_X15Y129_SLICE_X20Y129_BO6),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_CQ),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaeeeae)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_BLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_BQ),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a4b4b4b5a5a5a5a)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_ALUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I1(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_BQ),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I5(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y130_SLICE_X18Y130_AO6),
.Q(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hce3b0ace00000000)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X18Y130_CO5),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000008888)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_CLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I1(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777377708080808)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_BLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcd0101dccd1001)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_BO6),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_DQ),
.I5(CLBLM_R_X13Y130_SLICE_X18Y130_CO6),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.Q(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0b0e0f0f0f0f0f)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_CO6),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9d119d9da8a8a8a8)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.I4(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ff3737373f)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_CO5),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0033332121)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_ALUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_DO6),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y131_SLICE_X18Y131_AO6),
.Q(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y131_SLICE_X18Y131_BO6),
.Q(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0b0f0d0f)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.I1(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_CQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_DO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000011b099bb88)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_CLUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefa5450fefe5454)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_CO6),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I5(CLBLM_R_X13Y131_SLICE_X18Y131_CO6),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_BO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcced00330021)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_ALUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I5(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.Q(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555455ffffffff)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BQ),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_DO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000005040)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_CLUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_DQ),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_CO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55454555aababaaa)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_BLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I1(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_BQ),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.I5(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_BO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3330aaaa3330)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_A5Q),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00af00af00af00af)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I1(1'b1),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_DO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_CO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_BO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_ALUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_BQ),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I3(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_CQ),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_AO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_DO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_CO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_BO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_AO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000030)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_CQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_CO6),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_BQ),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_DO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fffffffffffffff)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_CQ),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_BQ),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_CO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_BLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_CO6),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_BQ),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I4(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_CQ),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_BO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c1e3c3c3c0f3c3c)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_ALUT (
.I0(CLBLM_R_X15Y129_SLICE_X20Y129_DO6),
.I1(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.I2(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I5(CLBLM_R_X15Y129_SLICE_X20Y129_CO6),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_AO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_DO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_CO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_BO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_AO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X15Y130_SLICE_X20Y130_AO6),
.Q(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_DO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_CO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_BO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcf000)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_DQ),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.I3(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.I4(CLBLM_R_X15Y129_SLICE_X20Y129_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_AO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X15Y130_SLICE_X21Y130_AO6),
.Q(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_DO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_CO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_BO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff3033fcfc3030)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I4(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_AO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X15Y132_SLICE_X20Y132_AO6),
.Q(CLBLM_R_X15Y132_SLICE_X20Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X20Y132_DO5),
.O6(CLBLM_R_X15Y132_SLICE_X20Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X20Y132_CO5),
.O6(CLBLM_R_X15Y132_SLICE_X20Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X20Y132_BO5),
.O6(CLBLM_R_X15Y132_SLICE_X20Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff400f4fff400f4)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X15Y132_SLICE_X20Y132_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X20Y132_AO5),
.O6(CLBLM_R_X15Y132_SLICE_X20Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X21Y132_DO5),
.O6(CLBLM_R_X15Y132_SLICE_X21Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X21Y132_CO5),
.O6(CLBLM_R_X15Y132_SLICE_X21Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X21Y132_BO5),
.O6(CLBLM_R_X15Y132_SLICE_X21Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X21Y132_AO5),
.O6(CLBLM_R_X15Y132_SLICE_X21Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y139_SLICE_X162Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y139_SLICE_X162Y139_DO5),
.O6(CLBLM_R_X103Y139_SLICE_X162Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y139_SLICE_X162Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y139_SLICE_X162Y139_CO5),
.O6(CLBLM_R_X103Y139_SLICE_X162Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y139_SLICE_X162Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y139_SLICE_X162Y139_BO5),
.O6(CLBLM_R_X103Y139_SLICE_X162Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y139_SLICE_X162Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y139_SLICE_X162Y139_AO5),
.O6(CLBLM_R_X103Y139_SLICE_X162Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y139_SLICE_X163Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y139_SLICE_X163Y139_DO5),
.O6(CLBLM_R_X103Y139_SLICE_X163Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y139_SLICE_X163Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y139_SLICE_X163Y139_CO5),
.O6(CLBLM_R_X103Y139_SLICE_X163Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y139_SLICE_X163Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y139_SLICE_X163Y139_BO5),
.O6(CLBLM_R_X103Y139_SLICE_X163Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00088880000)
  ) CLBLM_R_X103Y139_SLICE_X163Y139_ALUT (
.I0(RIOB33_X105Y139_IOB_X1Y140_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y137_IOB_X1Y138_I),
.I3(RIOB33_X105Y139_IOB_X1Y139_I),
.I4(RIOB33_X105Y141_IOB_X1Y141_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y139_SLICE_X163Y139_AO5),
.O6(CLBLM_R_X103Y139_SLICE_X163Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffccccffff)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffff00ffff)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffff0f0ffff)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X15Y132_SLICE_X20Y132_AQ),
.I3(CLBLM_R_X13Y122_SLICE_X19Y122_BQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_DO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_CO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_BO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_AO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_DO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_CO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_BO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffeeffee)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(1'b1),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_AO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffaaaaffff)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X0Y122_BO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X4Y128_SLICE_X5Y128_CO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_R_X11Y122_SLICE_X14Y122_A5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X4Y123_SLICE_X5Y123_CQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X4Y123_SLICE_X5Y123_DQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X10Y127_SLICE_X13Y127_D5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X4Y123_SLICE_X5Y123_D5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X11Y125_SLICE_X14Y125_C5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y128_SLICE_X2Y128_AQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X2Y131_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y130_SLICE_X2Y130_BQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X3Y128_SLICE_X2Y128_BQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y139_SLICE_X163Y139_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_R_X103Y139_SLICE_X163Y139_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X10Y153_SLICE_X13Y153_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X0Y123_AO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLL_L_X36Y127_SLICE_X54Y127_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X12Y129_SLICE_X16Y129_CO6),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X10Y153_SLICE_X13Y153_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X11Y137_SLICE_X14Y137_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X12Y129_SLICE_X16Y129_CO6),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y122_SLICE_X19Y122_BQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X15Y132_SLICE_X20Y132_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X103Y176_SLICE_X163Y176_AO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X103Y176_SLICE_X163Y176_AO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X15Y132_SLICE_X20Y132_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_AMUX = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_AMUX = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_BMUX = CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_AMUX = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B = CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D = CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A = CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B = CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C = CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D = CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_CMUX = CLBLL_L_X4Y123_SLICE_X5Y123_C5Q;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_DMUX = CLBLL_L_X4Y123_SLICE_X5Y123_D5Q;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_AMUX = CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_BMUX = CLBLL_L_X4Y124_SLICE_X4Y124_B5Q;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_CMUX = CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A = CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B = CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_CMUX = CLBLL_L_X4Y124_SLICE_X5Y124_CO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A = CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_BMUX = CLBLL_L_X4Y125_SLICE_X4Y125_B5Q;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_DMUX = CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A = CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_CMUX = CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_CMUX = CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A = CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B = CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_CMUX = CLBLL_L_X4Y127_SLICE_X4Y127_C5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A = CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_AMUX = CLBLL_L_X4Y127_SLICE_X5Y127_A5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_DMUX = CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B = CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C = CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D = CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_BMUX = CLBLL_L_X4Y128_SLICE_X4Y128_B5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_CMUX = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_DMUX = CLBLL_L_X4Y128_SLICE_X4Y128_D5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A = CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B = CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_AMUX = CLBLL_L_X4Y128_SLICE_X5Y128_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_BMUX = CLBLL_L_X4Y128_SLICE_X5Y128_BO5;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_CMUX = CLBLL_L_X4Y128_SLICE_X5Y128_CO5;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_DMUX = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A = CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_AMUX = CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_BMUX = CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B = CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CMUX = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_AMUX = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_BMUX = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_CMUX = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_AMUX = CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_CMUX = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B = CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_AMUX = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_AMUX = CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_BMUX = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B = CLBLL_L_X36Y127_SLICE_X54Y127_BO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C = CLBLL_L_X36Y127_SLICE_X54Y127_CO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D = CLBLL_L_X36Y127_SLICE_X54Y127_DO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A = CLBLL_L_X36Y127_SLICE_X55Y127_AO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B = CLBLL_L_X36Y127_SLICE_X55Y127_BO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C = CLBLL_L_X36Y127_SLICE_X55Y127_CO6;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D = CLBLL_L_X36Y127_SLICE_X55Y127_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_AMUX = CLBLM_L_X8Y121_SLICE_X10Y121_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_DMUX = CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_BMUX = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_DMUX = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A = CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_DMUX = CLBLM_L_X8Y122_SLICE_X11Y122_D5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_AMUX = CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_BMUX = CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A = CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B = CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CMUX = CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A = CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A = CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_DMUX = CLBLM_L_X8Y125_SLICE_X10Y125_D5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A = CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_AMUX = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_DMUX = CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_BMUX = CLBLM_L_X8Y126_SLICE_X10Y126_B5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CMUX = CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A = CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A = CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B = CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_CMUX = CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A = CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B = CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_CMUX = CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A = CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B = CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C = CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A = CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B = CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_BMUX = CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_AMUX = CLBLM_L_X8Y130_SLICE_X11Y130_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_AMUX = CLBLM_L_X8Y133_SLICE_X10Y133_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_DMUX = CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A = CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B = CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_AMUX = CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_BMUX = CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_BMUX = CLBLM_L_X10Y122_SLICE_X13Y122_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_CMUX = CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_AMUX = CLBLM_L_X10Y124_SLICE_X12Y124_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CMUX = CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_BMUX = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CMUX = CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A = CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_BMUX = CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A = CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_BMUX = CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_DMUX = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A = CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B = CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C = CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_AMUX = CLBLM_L_X10Y127_SLICE_X12Y127_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_BMUX = CLBLM_L_X10Y127_SLICE_X12Y127_B5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_DMUX = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A = CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_BMUX = CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_DMUX = CLBLM_L_X10Y127_SLICE_X13Y127_D5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_CMUX = CLBLM_L_X10Y128_SLICE_X12Y128_C5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_CMUX = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B = CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_CMUX = CLBLM_L_X10Y129_SLICE_X12Y129_C5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_DMUX = CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A = CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_AMUX = CLBLM_L_X10Y130_SLICE_X13Y130_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CMUX = CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CMUX = CLBLM_L_X10Y132_SLICE_X13Y132_C5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A = CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_BMUX = CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A = CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_BMUX = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_CMUX = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_AMUX = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A = CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B = CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C = CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B = CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C = CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D = CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_AMUX = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_BMUX = CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A = CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B = CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_AMUX = CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A = CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A = CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B = CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_AMUX = CLBLM_L_X12Y123_SLICE_X16Y123_A5Q;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_BMUX = CLBLM_L_X12Y123_SLICE_X16Y123_BO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_DMUX = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A = CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B = CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_AMUX = CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A = CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B = CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C = CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_CMUX = CLBLM_L_X12Y125_SLICE_X16Y125_C5Q;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A = CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B = CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D = CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_AMUX = CLBLM_L_X12Y125_SLICE_X17Y125_A5Q;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_BMUX = CLBLM_L_X12Y125_SLICE_X17Y125_B5Q;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_CMUX = CLBLM_L_X12Y125_SLICE_X17Y125_CO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_AMUX = CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_BMUX = CLBLM_L_X12Y126_SLICE_X16Y126_B5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_CMUX = CLBLM_L_X12Y126_SLICE_X16Y126_CO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A = CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B = CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_AMUX = CLBLM_L_X12Y127_SLICE_X16Y127_A5Q;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_BMUX = CLBLM_L_X12Y127_SLICE_X16Y127_BO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_DMUX = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A = CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C = CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D = CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A = CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B = CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D = CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_CMUX = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D = CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A = CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_AMUX = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_BMUX = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A = CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_BMUX = CLBLM_L_X12Y131_SLICE_X17Y131_BO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_CMUX = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_BMUX = CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_DMUX = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A = CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A = CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B = CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C = CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C = CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B = CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_AMUX = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A = CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C = CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_AMUX = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_AMUX = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B = CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_AMUX = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_DMUX = CLBLM_R_X3Y127_SLICE_X3Y127_DO5;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B = CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C = CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D = CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C = CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D = CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B = CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_CMUX = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A = CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C = CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_AMUX = CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_CMUX = CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_DMUX = CLBLM_R_X3Y130_SLICE_X2Y130_DO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D = CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_AMUX = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_BMUX = CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_AMUX = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CMUX = CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_BMUX = CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A = CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_AMUX = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_BMUX = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CMUX = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_DMUX = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A = CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_CMUX = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_AMUX = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_BMUX = CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A = CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B = CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C = CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A = CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B = CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C = CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_AMUX = CLBLM_R_X5Y123_SLICE_X7Y123_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_DMUX = CLBLM_R_X5Y123_SLICE_X7Y123_DO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A = CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_BMUX = CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A = CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_BMUX = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A = CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_BMUX = CLBLM_R_X5Y125_SLICE_X6Y125_B5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CMUX = CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_AMUX = CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AMUX = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_BMUX = CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_CMUX = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A = CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B = CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A = CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B = CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A = CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A = CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B = CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C = CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_AMUX = CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_AMUX = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_BMUX = CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_AMUX = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CMUX = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_DMUX = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A = CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B = CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_BMUX = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A = CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B = CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CMUX = CLBLM_R_X7Y124_SLICE_X8Y124_C5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_DMUX = CLBLM_R_X7Y124_SLICE_X8Y124_D5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A = CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B = CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_AMUX = CLBLM_R_X7Y124_SLICE_X9Y124_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_BMUX = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CMUX = CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_BMUX = CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CMUX = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_DMUX = CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CMUX = CLBLM_R_X7Y127_SLICE_X8Y127_C5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_DMUX = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_AMUX = CLBLM_R_X7Y127_SLICE_X9Y127_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A = CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B = CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C = CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_CMUX = CLBLM_R_X7Y128_SLICE_X8Y128_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A = CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_AMUX = CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CMUX = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A = CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_BMUX = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_AMUX = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_BMUX = CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_DMUX = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A = CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B = CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_AMUX = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_BMUX = CLBLM_R_X7Y139_SLICE_X9Y139_B5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CMUX = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_DMUX = CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A = CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_AMUX = CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_BMUX = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_AMUX = CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_BMUX = CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_AMUX = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_AMUX = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_CMUX = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_DMUX = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A = CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A = CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_BMUX = CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CMUX = CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A = CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_AMUX = CLBLM_R_X11Y126_SLICE_X14Y126_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_BMUX = CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CMUX = CLBLM_R_X11Y126_SLICE_X14Y126_C5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_DMUX = CLBLM_R_X11Y126_SLICE_X14Y126_D5Q;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A = CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A = CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_BMUX = CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_DMUX = CLBLM_R_X11Y127_SLICE_X14Y127_D5Q;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A = CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_AMUX = CLBLM_R_X11Y128_SLICE_X14Y128_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A = CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_AMUX = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_CMUX = CLBLM_R_X11Y128_SLICE_X15Y128_C5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_DMUX = CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A = CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_BMUX = CLBLM_R_X11Y129_SLICE_X14Y129_BO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B = CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_BMUX = CLBLM_R_X11Y130_SLICE_X14Y130_B5Q;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A = CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_AMUX = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_AMUX = CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_BMUX = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A = CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_AMUX = CLBLM_R_X11Y132_SLICE_X14Y132_A5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_CMUX = CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_AMUX = CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_BMUX = CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_AMUX = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_BMUX = CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_CMUX = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A = CLBLM_R_X13Y121_SLICE_X18Y121_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B = CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C = CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A = CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B = CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C = CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D = CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A = CLBLM_R_X13Y122_SLICE_X18Y122_AO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B = CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_AMUX = CLBLM_R_X13Y122_SLICE_X18Y122_AO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A = CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B = CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C = CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A = CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B = CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A = CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B = CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C = CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D = CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A = CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B = CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C = CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_AMUX = CLBLM_R_X13Y124_SLICE_X18Y124_A5Q;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_BMUX = CLBLM_R_X13Y124_SLICE_X18Y124_BO5;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A = CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B = CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D = CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A = CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C = CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D = CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_AMUX = CLBLM_R_X13Y125_SLICE_X18Y125_AO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_BMUX = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_CMUX = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A = CLBLM_R_X13Y125_SLICE_X19Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C = CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D = CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B = CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C = CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_CMUX = CLBLM_R_X13Y126_SLICE_X18Y126_CO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_DMUX = CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A = CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B = CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C = CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D = CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D = CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B = CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B = CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_CMUX = CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A = CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A = CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_BMUX = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_CMUX = CLBLM_R_X13Y130_SLICE_X18Y130_CO5;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D = CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_BMUX = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_CMUX = CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A = CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B = CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D = CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_CMUX = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B = CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C = CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D = CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D = CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B = CLBLM_R_X15Y128_SLICE_X20Y128_BO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A = CLBLM_R_X15Y128_SLICE_X21Y128_AO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D = CLBLM_R_X15Y128_SLICE_X21Y128_DO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A = CLBLM_R_X15Y129_SLICE_X20Y129_AO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B = CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C = CLBLM_R_X15Y129_SLICE_X20Y129_CO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D = CLBLM_R_X15Y129_SLICE_X20Y129_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A = CLBLM_R_X15Y129_SLICE_X21Y129_AO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C = CLBLM_R_X15Y129_SLICE_X21Y129_CO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A = CLBLM_R_X15Y130_SLICE_X20Y130_AO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B = CLBLM_R_X15Y130_SLICE_X20Y130_BO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C = CLBLM_R_X15Y130_SLICE_X20Y130_CO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D = CLBLM_R_X15Y130_SLICE_X20Y130_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A = CLBLM_R_X15Y130_SLICE_X21Y130_AO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B = CLBLM_R_X15Y130_SLICE_X21Y130_BO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C = CLBLM_R_X15Y130_SLICE_X21Y130_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D = CLBLM_R_X15Y130_SLICE_X21Y130_DO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A = CLBLM_R_X15Y132_SLICE_X20Y132_AO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B = CLBLM_R_X15Y132_SLICE_X20Y132_BO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C = CLBLM_R_X15Y132_SLICE_X20Y132_CO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D = CLBLM_R_X15Y132_SLICE_X20Y132_DO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A = CLBLM_R_X15Y132_SLICE_X21Y132_AO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B = CLBLM_R_X15Y132_SLICE_X21Y132_BO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C = CLBLM_R_X15Y132_SLICE_X21Y132_CO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D = CLBLM_R_X15Y132_SLICE_X21Y132_DO6;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_A = CLBLM_R_X103Y139_SLICE_X162Y139_AO6;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_B = CLBLM_R_X103Y139_SLICE_X162Y139_BO6;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_C = CLBLM_R_X103Y139_SLICE_X162Y139_CO6;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_D = CLBLM_R_X103Y139_SLICE_X162Y139_DO6;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_A = CLBLM_R_X103Y139_SLICE_X163Y139_AO6;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_B = CLBLM_R_X103Y139_SLICE_X163Y139_BO6;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_C = CLBLM_R_X103Y139_SLICE_X163Y139_CO6;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_D = CLBLM_R_X103Y139_SLICE_X163Y139_DO6;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_AMUX = CLBLM_R_X103Y139_SLICE_X163Y139_AO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_AMUX = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A = CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B = CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C = CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D = CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B = CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C = CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D = CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_AMUX = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A = CLBLM_R_X103Y176_SLICE_X162Y176_AO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B = CLBLM_R_X103Y176_SLICE_X162Y176_BO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C = CLBLM_R_X103Y176_SLICE_X162Y176_CO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D = CLBLM_R_X103Y176_SLICE_X162Y176_DO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B = CLBLM_R_X103Y176_SLICE_X163Y176_BO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C = CLBLM_R_X103Y176_SLICE_X163Y176_CO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D = CLBLM_R_X103Y176_SLICE_X163Y176_DO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X4Y123_SLICE_X5Y123_DQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X10Y127_SLICE_X13Y127_D5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X4Y123_SLICE_X5Y123_D5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y128_SLICE_X2Y128_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X3Y128_SLICE_X2Y128_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y139_SLICE_X163Y139_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_R_X103Y139_SLICE_X163Y139_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y130_SLICE_X2Y130_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y122_SLICE_X19Y122_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = CLBLM_R_X11Y130_SLICE_X15Y130_CQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A1 = CLBLM_R_X7Y139_SLICE_X9Y139_B5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A2 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A3 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A5 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_B5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B2 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B3 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B5 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A5 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A6 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C1 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B1 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B2 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B3 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B4 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B5 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B6 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C1 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C2 = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C4 = CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C5 = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C6 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D1 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D2 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D3 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D5 = CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D6 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A1 = CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A2 = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A3 = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A4 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A5 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A6 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B1 = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B2 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B3 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B4 = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B6 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C2 = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C3 = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C5 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C6 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D3 = CLBLM_L_X12Y125_SLICE_X16Y125_C5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D4 = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D5 = CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D4 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D6 = CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = CLBLM_L_X8Y129_SLICE_X10Y129_DQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = CLBLL_L_X4Y128_SLICE_X4Y128_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A1 = CLBLM_R_X7Y127_SLICE_X9Y127_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A3 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B3 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B5 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B6 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C3 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C4 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C5 = CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D1 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D2 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D3 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D6 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A2 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A5 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C1 = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C2 = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C3 = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C4 = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C5 = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C6 = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D1 = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D2 = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D4 = CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D6 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D6 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C4 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A1 = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A2 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A4 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A5 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A6 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B1 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B2 = CLBLM_R_X7Y130_SLICE_X8Y130_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C1 = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C2 = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C3 = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C4 = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C5 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C6 = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D2 = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D3 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D4 = CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D5 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D6 = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B1 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B2 = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B3 = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B5 = CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B6 = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C1 = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C2 = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C3 = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C4 = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C5 = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C6 = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D1 = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D3 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A1 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B1 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D4 = CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A1 = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A2 = CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A3 = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A4 = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A5 = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A6 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B1 = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B3 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B4 = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B5 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B6 = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C4 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C5 = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C6 = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D6 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D3 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D4 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C4 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C5 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C5 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A1 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A3 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A5 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C3 = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C4 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C5 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C6 = CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B2 = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A3 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B4 = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B1 = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B2 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B3 = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A1 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A2 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C1 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C2 = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C3 = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B3 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B4 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B5 = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B6 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D4 = CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D6 = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D2 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D3 = CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D4 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D5 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A2 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A4 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D2 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A6 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D3 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B2 = CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B3 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B4 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B5 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C2 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C3 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C4 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C5 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C6 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A2 = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A4 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_A1 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_A3 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_A4 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_A5 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_A6 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_B1 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_B2 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_B3 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_B4 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_B5 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_B6 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_C1 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_C2 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_C3 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_C4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_C5 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_D1 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_D2 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_D3 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_D4 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_D5 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X163Y139_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_A1 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_A2 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_A3 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_A4 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_A5 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_A6 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_B1 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_B2 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_B3 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_B4 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_B5 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_B6 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_C1 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_C2 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_C3 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_C4 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_C5 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_C6 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_D1 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_D2 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_D3 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_D4 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_D5 = 1'b1;
  assign CLBLM_R_X103Y139_SLICE_X162Y139_D6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A1 = CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A3 = CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A5 = CLBLL_L_X4Y126_SLICE_X4Y126_BQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A6 = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B4 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A1 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B5 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A5 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C6 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A1 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A2 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A3 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A4 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A5 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C5 = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B2 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B3 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B4 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B6 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C2 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C3 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C4 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C5 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D2 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D3 = CLBLM_L_X12Y121_SLICE_X17Y121_DQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D4 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A1 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A3 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A5 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B1 = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B2 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B3 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B5 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C1 = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C2 = CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C3 = CLBLM_L_X12Y123_SLICE_X16Y123_A5Q;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C4 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D1 = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D2 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D3 = CLBLM_L_X12Y126_SLICE_X16Y126_B5Q;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D4 = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D6 = CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A6 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A3 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A4 = CLBLL_L_X4Y128_SLICE_X4Y128_B5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_AX = CLBLM_R_X3Y127_SLICE_X3Y127_DO5;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B2 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B3 = CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B6 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C1 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C2 = CLBLM_R_X3Y127_SLICE_X3Y127_CQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C3 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C5 = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C6 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D2 = CLBLM_R_X3Y127_SLICE_X3Y127_CQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D4 = CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D5 = CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A1 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A3 = CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A6 = CLBLL_L_X4Y123_SLICE_X5Y123_DQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B1 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B2 = CLBLM_R_X3Y127_SLICE_X2Y127_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B3 = CLBLL_L_X4Y127_SLICE_X4Y127_DQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C1 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C2 = CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C3 = CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C5 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C6 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D3 = CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D4 = CLBLM_R_X3Y127_SLICE_X3Y127_CQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D6 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A2 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A3 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A4 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B1 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B2 = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B3 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B4 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B5 = CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B6 = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C2 = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C3 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C4 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C5 = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D1 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D2 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D6 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A1 = CLBLM_R_X5Y123_SLICE_X7Y123_A5Q;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A5 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A6 = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B2 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B3 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B4 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B5 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C3 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C4 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C5 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C6 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D1 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D2 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D4 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D5 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D6 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A2 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A3 = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A4 = CLBLM_R_X3Y128_SLICE_X2Y128_BQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A5 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A2 = CLBLM_R_X3Y128_SLICE_X2Y128_BQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A3 = CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A4 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A5 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A6 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B1 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B2 = CLBLM_R_X3Y128_SLICE_X2Y128_BQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B3 = CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B4 = CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A1 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A3 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A5 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B2 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B4 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B6 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C2 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C3 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C4 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C5 = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D2 = CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D4 = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D5 = CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D6 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A1 = CLBLM_R_X11Y128_SLICE_X14Y128_A5Q;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A2 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A5 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B1 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B2 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B3 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B4 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B5 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C3 = CLBLM_L_X12Y127_SLICE_X16Y127_DQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C2 = CLBLM_L_X12Y124_SLICE_X16Y124_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C3 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C4 = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C5 = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C6 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y139_SLICE_X163Y139_AO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D2 = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D3 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D4 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D5 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D6 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A1 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A3 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A4 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A6 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B1 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B2 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B3 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B4 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C1 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B1 = CLBLM_R_X11Y132_SLICE_X15Y132_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D1 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D2 = CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D3 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A3 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A4 = CLBLM_R_X3Y130_SLICE_X2Y130_DO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A5 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A6 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B1 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B2 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B5 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B6 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C1 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A3 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A4 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A6 = CLBLM_L_X12Y121_SLICE_X17Y121_DQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B1 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B2 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B5 = CLBLM_R_X11Y132_SLICE_X15Y132_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B6 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C2 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C4 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C5 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C6 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D1 = CLBLM_L_X12Y123_SLICE_X16Y123_A5Q;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D3 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D4 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D5 = CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D6 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A3 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A4 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A6 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_R_X103Y139_SLICE_X163Y139_AO5;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B2 = CLBLM_L_X12Y124_SLICE_X16Y124_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B3 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B4 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B5 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C2 = CLBLM_L_X12Y124_SLICE_X16Y124_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C4 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C6 = CLBLM_R_X11Y128_SLICE_X14Y128_A5Q;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D3 = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D2 = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D4 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D3 = CLBLM_L_X12Y124_SLICE_X16Y124_DQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D4 = CLBLM_L_X12Y124_SLICE_X16Y124_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A2 = CLBLM_R_X13Y128_SLICE_X19Y128_BQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A3 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A4 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A5 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A6 = CLBLM_R_X13Y128_SLICE_X18Y128_CQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A1 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C3 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C4 = CLBLL_L_X4Y126_SLICE_X4Y126_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C5 = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C4 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C5 = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A2 = CLBLM_R_X3Y128_SLICE_X2Y128_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A3 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A4 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A5 = CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A6 = CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_AX = CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B1 = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B2 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B5 = CLBLM_L_X10Y127_SLICE_X12Y127_A5Q;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B6 = CLBLM_R_X3Y130_SLICE_X2Y130_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C2 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C3 = CLBLM_R_X3Y130_SLICE_X2Y130_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C4 = CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C5 = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D1 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D2 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D3 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D4 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D5 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A1 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A3 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A4 = CLBLM_L_X12Y125_SLICE_X17Y125_DQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A5 = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D2 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_AX = CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D3 = CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B1 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B2 = CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B4 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B5 = CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D5 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_BX = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C1 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C4 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C5 = CLBLM_L_X12Y125_SLICE_X17Y125_B5Q;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D6 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D1 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D4 = CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D6 = CLBLM_L_X12Y125_SLICE_X17Y125_DQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A1 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A2 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A3 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A4 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A5 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B2 = CLBLM_L_X10Y130_SLICE_X13Y130_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B3 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B4 = CLBLM_R_X13Y125_SLICE_X19Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B5 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C1 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C2 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C3 = CLBLM_L_X12Y127_SLICE_X16Y127_A5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C4 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D1 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D2 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D3 = CLBLM_R_X13Y124_SLICE_X18Y124_BO5;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D4 = CLBLM_R_X13Y125_SLICE_X19Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D5 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D6 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y139_SLICE_X163Y139_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B3 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A2 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A3 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A4 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A5 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B4 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B3 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B4 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B5 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C2 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C3 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C4 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C5 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C6 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D2 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D3 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D4 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D5 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y130_SLICE_X2Y130_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A1 = CLBLM_R_X15Y129_SLICE_X20Y129_DO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A2 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A3 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A4 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A5 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A6 = CLBLM_R_X15Y129_SLICE_X20Y129_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B1 = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B2 = CLBLM_R_X13Y128_SLICE_X19Y128_BQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B3 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C4 = CLBLM_R_X11Y130_SLICE_X15Y130_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B4 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B5 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B6 = CLBLM_R_X13Y128_SLICE_X18Y128_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = CLBLM_R_X11Y130_SLICE_X14Y130_B5Q;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C5 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C2 = CLBLM_R_X13Y128_SLICE_X18Y128_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C3 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C4 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C5 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C6 = CLBLM_R_X13Y128_SLICE_X19Y128_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D2 = CLBLM_R_X13Y128_SLICE_X18Y128_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D3 = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D4 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D5 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D6 = CLBLM_R_X13Y128_SLICE_X19Y128_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A1 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A2 = CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A3 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A5 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B2 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C3 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C5 = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B3 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A2 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A3 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A5 = CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A6 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_AX = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B2 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B3 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B5 = CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C1 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C4 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C1 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D4 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D5 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D6 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A1 = CLBLM_R_X11Y126_SLICE_X14Y126_D5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A3 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C3 = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A6 = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B2 = CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B4 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B6 = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C2 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C3 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C4 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C6 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D1 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D2 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D4 = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D5 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D4 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A5 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A6 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_AX = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B1 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B3 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B5 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_BX = CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C1 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C2 = CLBLM_R_X13Y126_SLICE_X19Y126_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C5 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D2 = CLBLM_R_X11Y127_SLICE_X15Y127_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D3 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D4 = CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D5 = CLBLM_L_X12Y126_SLICE_X16Y126_B5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D6 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A3 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A4 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A5 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B6 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B4 = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B5 = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A1 = CLBLM_R_X11Y127_SLICE_X15Y127_DQ;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A2 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A3 = CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B6 = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A4 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A5 = CLBLM_R_X15Y129_SLICE_X20Y129_AO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B6 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A1 = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A2 = CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A3 = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A4 = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A5 = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A6 = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C4 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C5 = CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C1 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C2 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C5 = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A1 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B1 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C2 = CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C3 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D2 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D3 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D4 = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D6 = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A1 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A2 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A3 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A5 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B2 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B3 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C1 = CLBLL_L_X4Y127_SLICE_X4Y127_C5Q;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C2 = CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C3 = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D1 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D2 = CLBLM_L_X12Y127_SLICE_X17Y127_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D3 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D4 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D5 = CLBLM_R_X11Y127_SLICE_X15Y127_DQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A1 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A2 = CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A3 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_AX = CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B4 = CLBLM_R_X13Y127_SLICE_X18Y127_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B5 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C1 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C3 = CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C5 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D1 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D3 = CLBLM_L_X12Y127_SLICE_X16Y127_DQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D5 = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A3 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A4 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A5 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B5 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C5 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D5 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A1 = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A3 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A4 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A5 = CLBLM_L_X12Y130_SLICE_X16Y130_DQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A6 = CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B2 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B3 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B5 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B6 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C2 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C3 = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C4 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C5 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C6 = CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D1 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D2 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D3 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C6 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_R_X103Y139_SLICE_X163Y139_AO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A3 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A4 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A6 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B2 = CLBLM_L_X12Y128_SLICE_X17Y128_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B4 = CLBLM_R_X13Y128_SLICE_X18Y128_CQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C2 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D2 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A2 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A4 = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A5 = CLBLM_R_X13Y128_SLICE_X19Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A6 = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D2 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B1 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B2 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B3 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B5 = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C1 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C3 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C5 = CLBLM_L_X12Y127_SLICE_X16Y127_BO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D3 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D6 = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D4 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A1 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A2 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A4 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A5 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D5 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B1 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B2 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B4 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B5 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A1 = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A2 = CLBLM_R_X13Y122_SLICE_X19Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A3 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A5 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C1 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C2 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C3 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B2 = CLBLM_R_X13Y122_SLICE_X19Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B3 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B5 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B6 = CLBLM_L_X12Y123_SLICE_X16Y123_A5Q;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D1 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D2 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C1 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C2 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C3 = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C4 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C5 = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C6 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D4 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A1 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A3 = CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A5 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D1 = CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D2 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D3 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D4 = CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D5 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D6 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A6 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B1 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B2 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A1 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A2 = CLBLM_L_X12Y124_SLICE_X17Y124_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A3 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A5 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A6 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C1 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C2 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C3 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B2 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B5 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B6 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D1 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D2 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C1 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C2 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C3 = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C4 = CLBLM_R_X13Y122_SLICE_X18Y122_AO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C5 = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C6 = CLBLM_L_X12Y121_SLICE_X17Y121_CQ;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D4 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D5 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D1 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D2 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D3 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D4 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D5 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D6 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A1 = CLBLM_L_X10Y130_SLICE_X12Y130_DQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A2 = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A4 = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A5 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B2 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B3 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B4 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B5 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B6 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C4 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C2 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C3 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C4 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C5 = CLBLM_L_X12Y129_SLICE_X17Y129_CQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C6 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C5 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C6 = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D3 = CLBLM_L_X12Y129_SLICE_X17Y129_DQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D4 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D6 = CLBLM_R_X11Y127_SLICE_X15Y127_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A1 = CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A2 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A3 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A4 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A6 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B1 = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B2 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B6 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C1 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C2 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C3 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C4 = CLBLM_L_X12Y124_SLICE_X16Y124_DQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C5 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D3 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D6 = CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A3 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A5 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A6 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B2 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B3 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B4 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B5 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D6 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A2 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A3 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A6 = CLBLM_L_X12Y129_SLICE_X17Y129_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B2 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B3 = CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B6 = CLBLM_R_X11Y128_SLICE_X15Y128_BQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X4Y123_SLICE_X5Y123_D5Q;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C2 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C3 = CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C4 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C5 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D1 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D2 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D3 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D4 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D5 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D6 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A1 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A2 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A3 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A4 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_AX = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B1 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B2 = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B3 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B4 = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B5 = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B6 = CLBLM_L_X10Y130_SLICE_X13Y130_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C4 = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C2 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C3 = CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_SR = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A1 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A6 = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B1 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B2 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B4 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B5 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B6 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C2 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C3 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C5 = CLBLM_R_X7Y130_SLICE_X8Y130_CQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C6 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D1 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D5 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = CLBLM_L_X8Y122_SLICE_X11Y122_D5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A1 = CLBLM_R_X13Y123_SLICE_X19Y123_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A3 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A5 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A6 = CLBLM_R_X13Y128_SLICE_X19Y128_BQ;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D3 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D4 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A2 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A3 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A4 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A6 = CLBLM_R_X13Y124_SLICE_X18Y124_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_AX = CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B2 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B3 = CLBLM_L_X12Y124_SLICE_X16Y124_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B5 = CLBLM_R_X13Y124_SLICE_X18Y124_A5Q;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C2 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C3 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C5 = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C6 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D2 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D3 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D5 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D6 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C4 = CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C5 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A1 = CLBLM_L_X10Y131_SLICE_X13Y131_DQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A2 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A3 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A4 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A6 = CLBLM_L_X12Y131_SLICE_X16Y131_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B4 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B5 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B1 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C2 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B2 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B3 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B4 = CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B6 = CLBLM_R_X11Y128_SLICE_X15Y128_C5Q;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A1 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A3 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A6 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C2 = CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B1 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B3 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B4 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D2 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D3 = CLBLM_L_X12Y131_SLICE_X16Y131_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B6 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D5 = CLBLM_L_X12Y131_SLICE_X17Y131_BO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D6 = CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C1 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C2 = CLBLM_L_X8Y122_SLICE_X11Y122_D5Q;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C3 = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C4 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C6 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A1 = CLBLM_L_X12Y131_SLICE_X16Y131_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A6 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A3 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D1 = CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D2 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D3 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D4 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B5 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D6 = CLBLM_R_X7Y124_SLICE_X8Y124_D5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B1 = CLBLM_R_X11Y130_SLICE_X14Y130_DQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C2 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C3 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C4 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C5 = CLBLM_L_X12Y131_SLICE_X16Y131_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C6 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A1 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A2 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D1 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B2 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B3 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D1 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D5 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D6 = CLBLM_L_X12Y128_SLICE_X16Y128_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D3 = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D2 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D4 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C4 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D5 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D3 = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D4 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A2 = CLBLM_L_X12Y125_SLICE_X17Y125_CO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A3 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A5 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A6 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B2 = CLBLM_R_X13Y125_SLICE_X19Y125_BQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B3 = CLBLM_R_X13Y124_SLICE_X18Y124_A5Q;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B4 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B6 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D2 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A1 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A2 = CLBLM_L_X8Y121_SLICE_X10Y121_A5Q;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A3 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A4 = CLBLM_L_X12Y125_SLICE_X17Y125_A5Q;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_AX = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B1 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B2 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B3 = CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B4 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B5 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C1 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C2 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C3 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C4 = CLBLM_L_X12Y125_SLICE_X17Y125_BQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C5 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D3 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D4 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_SR = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A2 = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A4 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A5 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A6 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B1 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B2 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B4 = CLBLM_L_X12Y132_SLICE_X17Y132_CQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A1 = CLBLM_L_X10Y122_SLICE_X13Y122_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A2 = CLBLM_L_X12Y125_SLICE_X17Y125_DQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A3 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C4 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C5 = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C6 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C2 = CLBLM_L_X12Y132_SLICE_X17Y132_CQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B2 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B5 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C1 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C2 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C3 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A1 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A5 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A3 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A4 = CLBLM_L_X8Y130_SLICE_X11Y130_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D1 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B3 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B5 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D6 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B2 = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C2 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C5 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C6 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A3 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_AX = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B1 = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B5 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D2 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D5 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_BX = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D1 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C1 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C3 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C4 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C5 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C6 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D6 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D1 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D4 = CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D6 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A1 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A2 = CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A3 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A5 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A6 = CLBLM_R_X13Y125_SLICE_X18Y125_AO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B1 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B4 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B5 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B6 = CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X4Y123_SLICE_X5Y123_DQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C2 = CLBLM_R_X13Y126_SLICE_X19Y126_CQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C5 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C6 = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A3 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A4 = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A5 = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B2 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B3 = CLBLM_L_X12Y121_SLICE_X17Y121_DQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B4 = CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B5 = CLBLM_R_X13Y126_SLICE_X18Y126_CO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B6 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C1 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C3 = CLBLM_L_X12Y125_SLICE_X17Y125_A5Q;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C4 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C5 = CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D1 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D2 = CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D3 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D4 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D5 = CLBLM_L_X12Y125_SLICE_X17Y125_A5Q;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A2 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D6 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B2 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D2 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A1 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A2 = CLBLM_L_X12Y128_SLICE_X16Y128_DQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A4 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A5 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B1 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B2 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B3 = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B4 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B6 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C1 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C3 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D1 = CLBLM_L_X10Y130_SLICE_X13Y130_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D2 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D3 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D4 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D5 = CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D6 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = CLBLM_L_X12Y128_SLICE_X17Y128_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = CLBLM_L_X10Y129_SLICE_X12Y129_CQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A1 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A2 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A3 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A4 = CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A5 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A6 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B1 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B2 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B3 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B4 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B5 = CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B6 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A1 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A3 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A6 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B1 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C2 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C3 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D4 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D6 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_AX = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_AX = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B2 = 1'b1;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A1 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A3 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A6 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B1 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B3 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C4 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C5 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D2 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D4 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D6 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A1 = CLBLM_L_X10Y127_SLICE_X12Y127_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A2 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B1 = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B3 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B4 = CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B5 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B6 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C1 = CLBLM_R_X3Y125_SLICE_X3Y125_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C2 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C3 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C5 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_SR = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D1 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D3 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D4 = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A1 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A2 = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A4 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A5 = CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A6 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B1 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B2 = CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B3 = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B4 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B6 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D2 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C1 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C2 = CLBLM_R_X13Y128_SLICE_X19Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C3 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C4 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C5 = CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D5 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D1 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D2 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D3 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D5 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D6 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D6 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A2 = CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A3 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A4 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A5 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A6 = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B1 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B2 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B3 = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C1 = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C2 = CLBLM_R_X13Y128_SLICE_X18Y128_CQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C3 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C5 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C6 = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D1 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D2 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D3 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D5 = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_D5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C4 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A3 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C5 = CLBLM_L_X12Y132_SLICE_X17Y132_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A5 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B5 = CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X10Y127_SLICE_X13Y127_D5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B6 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B3 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A4 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A5 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A6 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D2 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D3 = CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B1 = CLBLM_L_X8Y124_SLICE_X11Y124_DQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B5 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D4 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C4 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C1 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C3 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C4 = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C5 = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C6 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C5 = CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D1 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D2 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D3 = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D4 = CLBLM_L_X10Y124_SLICE_X12Y124_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D5 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D6 = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A1 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A3 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A5 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B1 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B2 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B5 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C2 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C3 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C5 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D3 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D4 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D5 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D6 = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A1 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A2 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A3 = CLBLM_R_X13Y128_SLICE_X19Y128_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A4 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A5 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A6 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B1 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B2 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B3 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B4 = CLBLM_R_X13Y128_SLICE_X19Y128_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B5 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B6 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B6 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C1 = CLBLM_R_X13Y128_SLICE_X19Y128_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C2 = CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C3 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C4 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C5 = CLBLM_L_X12Y131_SLICE_X16Y131_CQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C6 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D1 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D2 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D3 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D4 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D5 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D6 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A1 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A2 = CLBLM_L_X12Y129_SLICE_X17Y129_CQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A3 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A5 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A6 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B1 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B2 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B3 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C4 = CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B4 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B6 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C5 = CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C1 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C2 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C3 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C4 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C5 = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C6 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D1 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D2 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D3 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D4 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D5 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D6 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A4 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A5 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A6 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B2 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B3 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B6 = CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C1 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C2 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A3 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A5 = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C3 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A6 = CLBLM_L_X10Y127_SLICE_X13Y127_D5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B1 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B2 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B3 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B4 = CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B5 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C5 = CLBLM_L_X10Y132_SLICE_X13Y132_C5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B6 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C2 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C3 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C4 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C5 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D1 = CLBLM_R_X11Y126_SLICE_X14Y126_C5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D3 = CLBLM_R_X7Y127_SLICE_X8Y127_C5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D5 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D6 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A1 = CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A3 = CLBLM_L_X12Y125_SLICE_X17Y125_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B2 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B3 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B4 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B5 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C2 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C5 = CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C6 = CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D3 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y130_SLICE_X2Y130_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D3 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D4 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D6 = CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D6 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A1 = CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A2 = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A3 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A5 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B1 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B2 = CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B3 = CLBLM_R_X13Y130_SLICE_X18Y130_CO5;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B4 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A1 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A3 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A6 = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C2 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C3 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D1 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D3 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D4 = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A3 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A4 = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_DQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A6 = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B1 = CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B2 = CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B3 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A2 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A3 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A5 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C1 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C2 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C3 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B2 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B3 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B5 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D1 = CLBLM_R_X13Y130_SLICE_X18Y130_CO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D2 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C3 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D3 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D5 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D6 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D1 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D3 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D5 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A2 = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A3 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A4 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A2 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A5 = CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C6 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A4 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A5 = CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A6 = CLBLM_L_X10Y128_SLICE_X12Y128_C5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_AX = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D4 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B5 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C6 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C2 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C4 = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B2 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B1 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B5 = CLBLM_R_X5Y123_SLICE_X7Y123_DO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D1 = CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D2 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D5 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C2 = CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C4 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D3 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D5 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A2 = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A3 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A4 = CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B1 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B2 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B3 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B4 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B5 = CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B6 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A3 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A5 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C1 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C2 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B2 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B3 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B4 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B5 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D1 = CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C1 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C2 = CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C4 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C5 = CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C6 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D3 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A1 = CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A3 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A4 = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A5 = CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A6 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D2 = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C3 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D3 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D4 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D5 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D6 = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C4 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B2 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A3 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A4 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A5 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C1 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C2 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C3 = CLBLM_L_X12Y131_SLICE_X16Y131_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B1 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B3 = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B4 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B5 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B6 = CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D1 = CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D2 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_D5Q;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C2 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C4 = CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C5 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C6 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D3 = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D4 = CLBLM_L_X12Y129_SLICE_X17Y129_CQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D5 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D6 = CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D1 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D2 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D3 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D4 = CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D5 = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D6 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A4 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A5 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B4 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B5 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B6 = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C1 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C3 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C4 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C5 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D4 = CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A4 = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A5 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B1 = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B4 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A1 = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A2 = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C5 = CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C1 = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B1 = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B5 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C1 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C2 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C4 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C5 = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D2 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D5 = CLBLM_R_X5Y123_SLICE_X7Y123_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D6 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D5 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A1 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A2 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A5 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A6 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B1 = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B3 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B4 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B5 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B6 = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C1 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C2 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C3 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C5 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D6 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A1 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D1 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D4 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D6 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B5 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A3 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A4 = CLBLM_R_X11Y126_SLICE_X14Y126_D5Q;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A5 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B2 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B3 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B4 = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A5 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C3 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C4 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C5 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D1 = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D2 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D4 = CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B2 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B4 = CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B5 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B6 = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_BX = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C3 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A1 = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C4 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A4 = CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A6 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C5 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A4 = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A5 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A1 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B1 = CLBLL_L_X4Y125_SLICE_X4Y125_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B4 = CLBLM_R_X3Y125_SLICE_X3Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B5 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D1 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D2 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D3 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D4 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D5 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D1 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A2 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A3 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A6 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D1 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B1 = CLBLM_L_X12Y129_SLICE_X17Y129_DQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B2 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B4 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A3 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A4 = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A5 = CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B6 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B2 = CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_CO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B4 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B5 = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A3 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C1 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C2 = CLBLM_R_X5Y123_SLICE_X7Y123_A5Q;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C3 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C5 = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D2 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D3 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D4 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D4 = CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D5 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D6 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C6 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B5 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_A5Q;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A2 = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A4 = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A5 = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A6 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D2 = CLBLM_R_X13Y128_SLICE_X18Y128_DQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B1 = CLBLM_L_X12Y123_SLICE_X16Y123_BO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B2 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B3 = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B4 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B5 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B6 = CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C3 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C1 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C2 = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C4 = CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C5 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C6 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D5 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D6 = CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y128_SLICE_X2Y128_AQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D1 = CLBLM_L_X8Y122_SLICE_X11Y122_D5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D2 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D3 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D4 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D5 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A2 = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A3 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A5 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B1 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B2 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B4 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B5 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C1 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C2 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C3 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C4 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C5 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C6 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_D5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D5 = CLBLM_L_X12Y126_SLICE_X16Y126_B5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D6 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A4 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C4 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C5 = CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C6 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D4 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B3 = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D5 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B4 = CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B5 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B6 = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A1 = CLBLL_L_X4Y124_SLICE_X4Y124_B5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A3 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B1 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B2 = CLBLL_L_X4Y126_SLICE_X4Y126_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B4 = CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B5 = CLBLM_L_X12Y124_SLICE_X17Y124_CQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B6 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C1 = CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C2 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C3 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C4 = CLBLM_R_X7Y128_SLICE_X8Y128_C5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_AX = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = CLBLM_L_X8Y124_SLICE_X11Y124_DQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = CLBLM_L_X10Y130_SLICE_X13Y130_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D3 = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D5 = CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = CLBLM_L_X12Y131_SLICE_X16Y131_DQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D5 = CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = CLBLM_R_X11Y130_SLICE_X15Y130_BQ;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A2 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A3 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A5 = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B2 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B3 = CLBLM_R_X5Y125_SLICE_X6Y125_B5Q;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B6 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C1 = CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C2 = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C4 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C5 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C6 = CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = CLBLM_R_X11Y130_SLICE_X15Y130_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D2 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D3 = CLBLL_L_X4Y128_SLICE_X5Y128_BO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D4 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D6 = CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B1 = CLBLM_R_X3Y128_SLICE_X2Y128_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B2 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B3 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A2 = CLBLM_R_X13Y123_SLICE_X18Y123_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A3 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A5 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B5 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B1 = CLBLM_L_X12Y125_SLICE_X16Y125_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B3 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C4 = CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B5 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B6 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C5 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C1 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C2 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C4 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C5 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C6 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D2 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D6 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A2 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A3 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A5 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C4 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C5 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B4 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B5 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C5 = CLBLM_L_X12Y126_SLICE_X16Y126_B5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C6 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D3 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D2 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D3 = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D4 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D5 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D5 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A1 = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A3 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A4 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B2 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B4 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C1 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C3 = CLBLL_L_X4Y127_SLICE_X4Y127_DQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C4 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = CLBLM_L_X12Y131_SLICE_X16Y131_DQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D1 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D3 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A4 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A5 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B4 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C3 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C4 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C5 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C6 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = CLBLM_L_X10Y131_SLICE_X13Y131_DQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A1 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A3 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D1 = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A5 = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D2 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D4 = CLBLM_L_X8Y122_SLICE_X11Y122_D5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D6 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A6 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_AX = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A2 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A3 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A6 = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_AX = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B2 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C2 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C5 = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C6 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D3 = CLBLM_R_X5Y125_SLICE_X6Y125_B5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D4 = CLBLL_L_X4Y127_SLICE_X5Y127_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D2 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D3 = CLBLM_L_X8Y121_SLICE_X10Y121_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D4 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A1 = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A2 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A3 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A5 = CLBLM_L_X8Y125_SLICE_X10Y125_D5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B4 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C2 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C4 = CLBLM_L_X12Y124_SLICE_X16Y124_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C5 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D2 = CLBLM_R_X13Y127_SLICE_X18Y127_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D3 = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D4 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D5 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A1 = CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A5 = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A6 = CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B1 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B2 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B5 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C1 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C5 = CLBLM_R_X11Y126_SLICE_X14Y126_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D2 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D4 = CLBLM_R_X13Y127_SLICE_X18Y127_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D5 = CLBLM_L_X10Y128_SLICE_X12Y128_DQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D6 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A1 = CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A2 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A3 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A4 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A6 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B3 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B5 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C2 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C3 = CLBLL_L_X4Y124_SLICE_X4Y124_B5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C4 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C5 = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = CLBLM_L_X10Y130_SLICE_X13Y130_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = CLBLM_R_X11Y128_SLICE_X15Y128_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D1 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D2 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A3 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A4 = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A5 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B2 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = CLBLM_L_X10Y130_SLICE_X13Y130_DQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B3 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B6 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C2 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C6 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A3 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A5 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_AX = CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B1 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B2 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B5 = CLBLL_L_X4Y128_SLICE_X5Y128_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C4 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D1 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D2 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D3 = CLBLL_L_X4Y128_SLICE_X4Y128_B5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D4 = CLBLL_L_X4Y127_SLICE_X5Y127_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D5 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D6 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C1 = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C6 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D3 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D4 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D5 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A1 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A2 = CLBLM_L_X12Y126_SLICE_X16Y126_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A4 = CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A6 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B1 = CLBLM_R_X13Y126_SLICE_X19Y126_CQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B2 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B4 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B6 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C3 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C5 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C6 = CLBLM_L_X10Y124_SLICE_X12Y124_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D2 = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D3 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D4 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D5 = CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A3 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A4 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_AX = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B2 = CLBLM_L_X10Y124_SLICE_X12Y124_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B4 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C2 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C4 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C5 = CLBLM_R_X11Y127_SLICE_X15Y127_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D1 = CLBLM_R_X11Y126_SLICE_X14Y126_C5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D2 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D3 = CLBLM_L_X10Y132_SLICE_X13Y132_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D6 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A3 = CLBLM_R_X3Y127_SLICE_X3Y127_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A4 = CLBLL_L_X4Y128_SLICE_X4Y128_DQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A6 = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_AX = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B1 = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B2 = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B3 = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B4 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B5 = CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B6 = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C1 = CLBLM_R_X3Y127_SLICE_X2Y127_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C2 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C3 = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C4 = CLBLL_L_X4Y125_SLICE_X4Y125_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A2 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A4 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D5 = CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D6 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A6 = CLBLM_L_X8Y131_SLICE_X10Y131_DQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B2 = CLBLM_R_X11Y126_SLICE_X14Y126_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B4 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A2 = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A3 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C1 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C2 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B1 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B2 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B3 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B4 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B5 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C1 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C2 = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C3 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C4 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B1 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D4 = CLBLM_L_X8Y124_SLICE_X11Y124_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C1 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C4 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A1 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A2 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A4 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A5 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D1 = CLBLL_L_X4Y127_SLICE_X5Y127_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D2 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D5 = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B1 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B3 = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B4 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B5 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_D5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C6 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D1 = CLBLM_L_X8Y121_SLICE_X10Y121_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D3 = CLBLM_L_X12Y128_SLICE_X17Y128_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D4 = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D5 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D6 = CLBLM_L_X8Y125_SLICE_X10Y125_D5Q;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A3 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A4 = CLBLM_R_X11Y128_SLICE_X15Y128_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A5 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A6 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B2 = CLBLM_R_X11Y127_SLICE_X15Y127_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B5 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B6 = CLBLM_R_X11Y127_SLICE_X14Y127_D5Q;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C2 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C3 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C4 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C5 = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D1 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D3 = CLBLM_R_X11Y127_SLICE_X15Y127_DQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D5 = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A1 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A2 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A3 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B1 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B2 = CLBLM_L_X12Y127_SLICE_X16Y127_DQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B3 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C2 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C3 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C5 = CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C6 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B2 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D2 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D3 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D4 = CLBLM_L_X8Y126_SLICE_X10Y126_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D6 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A3 = CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A4 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A5 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A6 = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C2 = CLBLL_L_X4Y125_SLICE_X4Y125_CQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C3 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B1 = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B2 = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B3 = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B4 = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B5 = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B6 = CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C1 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C3 = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C4 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C5 = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C6 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C6 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D2 = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D3 = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D4 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D5 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D6 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A2 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A5 = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A6 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B1 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B2 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B3 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B5 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B6 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A3 = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A4 = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C2 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C3 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C4 = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A5 = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A6 = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B2 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B3 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B4 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B5 = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B6 = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C2 = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C3 = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C4 = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C5 = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C6 = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D3 = CLBLM_L_X8Y124_SLICE_X11Y124_DQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D4 = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A2 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D2 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D4 = CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D5 = CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D6 = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A5 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A6 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B1 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B2 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B4 = CLBLL_L_X4Y128_SLICE_X4Y128_D5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C1 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C2 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C4 = CLBLM_L_X12Y123_SLICE_X17Y123_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C4 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C5 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D2 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D3 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D5 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C6 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A3 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A6 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_AX = CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B2 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B5 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B6 = CLBLM_R_X11Y128_SLICE_X15Y128_BQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C1 = CLBLM_R_X5Y123_SLICE_X7Y123_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C3 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D3 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D5 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D3 = CLBLM_L_X10Y130_SLICE_X12Y130_DQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D4 = CLBLM_L_X10Y130_SLICE_X13Y130_CQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D5 = CLBLM_R_X11Y130_SLICE_X14Y130_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A1 = CLBLM_R_X11Y127_SLICE_X14Y127_D5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A2 = CLBLM_R_X11Y128_SLICE_X14Y128_DQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_AX = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B1 = CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B2 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B3 = CLBLM_R_X11Y128_SLICE_X14Y128_DQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A1 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C1 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C3 = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C5 = CLBLM_L_X10Y128_SLICE_X12Y128_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D2 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D3 = CLBLM_R_X11Y128_SLICE_X14Y128_DQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D5 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A2 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A3 = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A4 = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A5 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A6 = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B1 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B2 = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B3 = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B4 = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B5 = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B6 = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C2 = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C3 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C5 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C6 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B6 = CLBLM_L_X10Y130_SLICE_X13Y130_A5Q;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D1 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D2 = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D3 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D4 = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D6 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A1 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A2 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D2 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D3 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A1 = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A2 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A3 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A4 = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A5 = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A6 = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B2 = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B3 = CLBLL_L_X4Y128_SLICE_X5Y128_CO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B4 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B5 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C3 = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C4 = CLBLM_L_X10Y128_SLICE_X12Y128_DQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C2 = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C3 = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C6 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D3 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D5 = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D2 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D3 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D5 = CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D6 = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A4 = CLBLM_R_X13Y125_SLICE_X19Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A5 = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B2 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B4 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B5 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B6 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C2 = CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C4 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C5 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D1 = CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D4 = CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D5 = CLBLM_L_X8Y125_SLICE_X10Y125_D5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B2 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D5 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A5 = CLBLM_L_X12Y127_SLICE_X16Y127_A5Q;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B2 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B3 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B5 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B6 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B6 = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C1 = CLBLM_R_X11Y130_SLICE_X15Y130_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C2 = CLBLM_R_X11Y130_SLICE_X14Y130_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C3 = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C4 = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C5 = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C6 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D2 = CLBLM_L_X12Y128_SLICE_X16Y128_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D3 = CLBLM_R_X11Y130_SLICE_X15Y130_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D4 = CLBLM_R_X11Y129_SLICE_X14Y129_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D5 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D6 = CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A2 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A3 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A4 = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C3 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B1 = CLBLM_R_X11Y130_SLICE_X14Y130_DQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B2 = CLBLM_R_X11Y130_SLICE_X14Y130_B5Q;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B5 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C4 = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C5 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C1 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C2 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C3 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C5 = CLBLM_R_X11Y129_SLICE_X14Y129_BO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C6 = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D2 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D3 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D4 = CLBLM_R_X11Y127_SLICE_X14Y127_CQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D5 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D6 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A1 = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A2 = CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A3 = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A4 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A6 = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B1 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B2 = CLBLM_R_X3Y127_SLICE_X2Y127_DQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B3 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B4 = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B5 = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B6 = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C1 = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C2 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C3 = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C4 = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C5 = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C6 = CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D1 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D2 = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A2 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A3 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A4 = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A6 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B1 = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B2 = CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B3 = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B5 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B6 = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B4 = CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B5 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C2 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C3 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C4 = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C5 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C6 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D1 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D2 = CLBLM_R_X7Y127_SLICE_X9Y127_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D6 = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D2 = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A4 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A6 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B1 = CLBLM_L_X8Y126_SLICE_X10Y126_B5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B2 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B5 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C1 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C2 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C3 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D1 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D2 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D3 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D4 = CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D5 = CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C4 = CLBLM_L_X10Y130_SLICE_X13Y130_CQ;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A1 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A3 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A4 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A5 = CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A6 = CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y122_SLICE_X19Y122_BQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_AX = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B4 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B5 = CLBLM_L_X12Y126_SLICE_X16Y126_CO5;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B6 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = CLBLL_L_X4Y123_SLICE_X5Y123_C5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C2 = CLBLM_R_X11Y130_SLICE_X15Y130_CQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C3 = CLBLM_L_X10Y132_SLICE_X13Y132_CQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D3 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D4 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A2 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A3 = CLBLM_L_X12Y129_SLICE_X17Y129_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B1 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C3 = CLBLM_L_X8Y129_SLICE_X10Y129_DQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D3 = CLBLM_R_X11Y130_SLICE_X14Y130_DQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D4 = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D5 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C1 = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C2 = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C4 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C5 = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C6 = CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D4 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D5 = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D6 = CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A5 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A2 = CLBLM_L_X8Y126_SLICE_X10Y126_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B2 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B4 = CLBLM_L_X10Y128_SLICE_X12Y128_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B5 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B6 = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C3 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C4 = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C5 = CLBLM_L_X10Y129_SLICE_X12Y129_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C4 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D1 = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D2 = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D6 = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D4 = CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A2 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A4 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A5 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A6 = CLBLM_L_X12Y128_SLICE_X17Y128_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B4 = CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B5 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C1 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C2 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C4 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D1 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D2 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D5 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D6 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = CLBLM_L_X12Y124_SLICE_X16Y124_DQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = CLBLM_R_X11Y132_SLICE_X15Y132_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_AX = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = CLBLM_L_X12Y126_SLICE_X17Y126_CQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_BX = CLBLM_R_X7Y127_SLICE_X9Y127_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = CLBLM_L_X10Y130_SLICE_X13Y130_DQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_CQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_SR = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B1 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B2 = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B4 = CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B5 = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B6 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C2 = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C5 = CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D1 = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D2 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D3 = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D4 = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D5 = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D6 = CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A3 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B3 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D4 = CLBLM_R_X7Y127_SLICE_X8Y127_C5Q;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A1 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A4 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A5 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B2 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B3 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B4 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B5 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C2 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C4 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C6 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D1 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D2 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D3 = CLBLM_L_X8Y128_SLICE_X10Y128_DQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A1 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A2 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A4 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A6 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B1 = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B2 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B4 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B5 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B6 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C1 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C2 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C3 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D6 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A1 = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A2 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A3 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A4 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_AX = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B2 = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B3 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B4 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C2 = CLBLM_L_X10Y130_SLICE_X13Y130_DQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = CLBLL_L_X4Y125_SLICE_X4Y125_B5Q;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D4 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D6 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X3Y128_SLICE_X2Y128_BQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A2 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A3 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A5 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A6 = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B1 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B5 = CLBLM_L_X8Y124_SLICE_X11Y124_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B6 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C2 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C3 = CLBLM_L_X10Y130_SLICE_X12Y130_DQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C5 = CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C6 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D1 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D3 = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D4 = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A2 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A5 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A6 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B2 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B5 = CLBLM_R_X11Y130_SLICE_X15Y130_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B6 = CLBLL_L_X4Y128_SLICE_X4Y128_DQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C1 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C2 = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C3 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C5 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D3 = CLBLM_L_X8Y129_SLICE_X10Y129_DQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D6 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A3 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A4 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A5 = CLBLM_L_X10Y130_SLICE_X13Y130_A5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B1 = CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B2 = CLBLM_L_X12Y132_SLICE_X17Y132_CQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B3 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D1 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B4 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B5 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A3 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C1 = CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C2 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C3 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B1 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B3 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B4 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D1 = CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D2 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C1 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C2 = CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C3 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C5 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C6 = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D3 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D4 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A1 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A2 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A4 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A5 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D1 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D4 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D5 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D6 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_AX = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B1 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B2 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B3 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B4 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A2 = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A4 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C1 = CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C2 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C3 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B2 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B5 = CLBLM_R_X7Y128_SLICE_X8Y128_C5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C3 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C4 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C5 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C6 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D4 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_SR = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D1 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D3 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D4 = CLBLM_L_X12Y125_SLICE_X17Y125_B5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D5 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D6 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A1 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B1 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = CLBLM_L_X12Y130_SLICE_X16Y130_DQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B4 = CLBLM_L_X12Y125_SLICE_X17Y125_B5Q;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B5 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A6 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B1 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B2 = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B3 = CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B4 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B5 = CLBLM_L_X12Y132_SLICE_X17Y132_CQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B6 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A1 = CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A3 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_AX = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B1 = CLBLM_R_X7Y124_SLICE_X8Y124_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B2 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B3 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C4 = CLBLM_R_X11Y130_SLICE_X15Y130_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_BX = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C5 = CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C1 = CLBLM_L_X10Y128_SLICE_X12Y128_C5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C4 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C5 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D4 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A6 = CLBLM_R_X11Y132_SLICE_X14Y132_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D1 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D2 = CLBLM_L_X8Y121_SLICE_X10Y121_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D4 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D5 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D6 = CLBLM_R_X3Y125_SLICE_X3Y125_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B2 = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B4 = CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B5 = CLBLM_L_X10Y130_SLICE_X13Y130_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A4 = CLBLM_R_X11Y125_SLICE_X15Y125_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A5 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C1 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C2 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B3 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B4 = CLBLM_L_X8Y124_SLICE_X11Y124_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C1 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C5 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D4 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D1 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D2 = CLBLM_R_X7Y124_SLICE_X9Y124_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D6 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A3 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A4 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = CLBLM_L_X10Y130_SLICE_X12Y130_DQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = CLBLL_L_X4Y128_SLICE_X4Y128_D5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = CLBLM_L_X8Y131_SLICE_X10Y131_DQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C4 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B5 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B6 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = CLBLM_L_X8Y126_SLICE_X10Y126_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D5 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X4Y123_SLICE_X5Y123_CQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X4Y123_SLICE_X5Y123_DQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X10Y127_SLICE_X13Y127_D5Q;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A1 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A2 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A3 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A4 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A6 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B1 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B2 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B5 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B6 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C4 = CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C5 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C6 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D1 = CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D3 = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D5 = CLBLM_L_X8Y131_SLICE_X10Y131_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D6 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A3 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A5 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A6 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B1 = CLBLM_R_X11Y127_SLICE_X14Y127_DQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B2 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B3 = CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C1 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C2 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C3 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C4 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D1 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D3 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D5 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A1 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A2 = CLBLM_L_X8Y126_SLICE_X10Y126_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A4 = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A5 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B1 = CLBLM_L_X10Y127_SLICE_X12Y127_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B5 = CLBLM_L_X10Y128_SLICE_X12Y128_C5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C1 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C2 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C4 = CLBLL_L_X4Y123_SLICE_X5Y123_C5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C5 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D1 = CLBLM_R_X11Y128_SLICE_X15Y128_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D2 = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D3 = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D4 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D6 = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = CLBLM_L_X10Y129_SLICE_X12Y129_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_AX = CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A3 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A4 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A2 = CLBLM_L_X12Y125_SLICE_X17Y125_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A3 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A6 = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_AX = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B1 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B2 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B4 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C1 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C3 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C5 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C6 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A2 = CLBLM_R_X11Y132_SLICE_X14Y132_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A5 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D2 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D3 = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D4 = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D6 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A2 = CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A4 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B2 = CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B3 = CLBLM_L_X12Y125_SLICE_X16Y125_C5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B4 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B5 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B6 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C1 = CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C4 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C5 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D2 = CLBLM_L_X10Y127_SLICE_X12Y127_B5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D4 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D5 = CLBLM_L_X10Y128_SLICE_X12Y128_C5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D6 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C4 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D5 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D6 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B5 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X4Y123_SLICE_X5Y123_D5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A2 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A3 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B2 = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B5 = CLBLM_L_X8Y124_SLICE_X11Y124_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C1 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C2 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C4 = CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C6 = CLBLM_L_X12Y126_SLICE_X17Y126_BQ;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D2 = CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D3 = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D4 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A3 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A4 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A6 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B2 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B6 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C1 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C2 = CLBLM_L_X10Y132_SLICE_X13Y132_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B2 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C4 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C5 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B3 = CLBLL_L_X4Y127_SLICE_X4Y127_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D2 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B5 = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D3 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D4 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D6 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B6 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C1 = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C2 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C3 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C6 = CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D5 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = CLBLM_R_X15Y132_SLICE_X20Y132_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = CLBLM_R_X13Y122_SLICE_X19Y122_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y128_SLICE_X2Y128_AQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = CLBLM_L_X8Y128_SLICE_X10Y128_DQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A2 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A3 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A4 = CLBLM_L_X8Y126_SLICE_X10Y126_BQ;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_A6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C3 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B1 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B2 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B3 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B4 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B5 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_B6 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C1 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C2 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C3 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C4 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C5 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_C6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D1 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D2 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D3 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D4 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D5 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X54Y127_D6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C5 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A1 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A2 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A3 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A4 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A5 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B1 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B2 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B3 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B4 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B5 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_B6 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C1 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C2 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C3 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C4 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C5 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_C6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D1 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D2 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D3 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D4 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D5 = 1'b1;
  assign CLBLL_L_X36Y127_SLICE_X55Y127_D6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = CLBLM_L_X12Y129_SLICE_X17Y129_DQ;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A4 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B1 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B4 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C1 = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C2 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C3 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C4 = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C5 = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C6 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D2 = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D5 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A2 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A4 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A6 = CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B1 = CLBLM_R_X11Y126_SLICE_X15Y126_DQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C1 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C2 = CLBLM_R_X7Y130_SLICE_X8Y130_CQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D1 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D3 = CLBLM_R_X7Y130_SLICE_X8Y130_DQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D5 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = CLBLM_L_X10Y131_SLICE_X13Y131_DQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C2 = CLBLM_L_X10Y129_SLICE_X12Y129_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C3 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D3 = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D5 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A2 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A4 = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A5 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B2 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B3 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y122_SLICE_X19Y122_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B4 = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = CLBLM_L_X8Y130_SLICE_X11Y130_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A1 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A3 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B1 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B2 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B4 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = CLBLM_R_X11Y125_SLICE_X15Y125_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B4 = CLBLM_L_X10Y128_SLICE_X12Y128_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A1 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A2 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A3 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A4 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A5 = CLBLM_R_X3Y130_SLICE_X2Y130_BQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A6 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B2 = CLBLM_R_X3Y131_SLICE_X2Y131_A5Q;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B6 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A1 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A4 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A5 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A6 = CLBLM_R_X7Y139_SLICE_X9Y139_B5Q;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D6 = 1'b1;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A1 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A2 = CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A3 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A5 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A2 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A5 = CLBLM_R_X11Y122_SLICE_X14Y122_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C2 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_AX = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B2 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B4 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B5 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B6 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C1 = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C2 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C6 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D4 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A3 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D3 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D4 = CLBLM_R_X5Y123_SLICE_X7Y123_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D5 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A6 = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A1 = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A2 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A3 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B1 = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B2 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B6 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D2 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C1 = CLBLL_L_X4Y123_SLICE_X5Y123_D5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C5 = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D4 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D2 = CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D4 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D6 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C5 = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C5 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C3 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C4 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_B5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CE = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A4 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A5 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A6 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B1 = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B3 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B4 = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B5 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B6 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C2 = CLBLL_L_X4Y128_SLICE_X4Y128_D5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C3 = CLBLM_R_X5Y125_SLICE_X6Y125_B5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C5 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C6 = CLBLM_L_X8Y130_SLICE_X11Y130_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D2 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D4 = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D5 = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D6 = CLBLM_L_X8Y130_SLICE_X11Y130_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A2 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A5 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A6 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C5 = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B2 = CLBLM_R_X3Y127_SLICE_X2Y127_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B3 = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B4 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B5 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C6 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C1 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C2 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C4 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D1 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D3 = CLBLM_R_X3Y128_SLICE_X2Y128_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D4 = CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D5 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D6 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = CLBLM_L_X10Y130_SLICE_X13Y130_DQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLL_L_X36Y127_SLICE_X54Y127_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = CLBLM_L_X10Y133_SLICE_X13Y133_B5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = CLBLL_L_X4Y128_SLICE_X5Y128_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = CLBLM_L_X12Y131_SLICE_X16Y131_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A1 = CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A2 = CLBLM_R_X5Y125_SLICE_X6Y125_B5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A3 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A4 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A5 = CLBLL_L_X4Y123_SLICE_X5Y123_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B1 = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B2 = CLBLM_R_X11Y128_SLICE_X15Y128_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B3 = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B4 = CLBLM_L_X8Y130_SLICE_X11Y130_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B5 = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C2 = CLBLM_R_X11Y128_SLICE_X15Y128_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C3 = CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C4 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C6 = CLBLL_L_X4Y128_SLICE_X4Y128_D5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X3Y128_SLICE_X2Y128_BQ;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D2 = CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D3 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D4 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D5 = CLBLL_L_X4Y123_SLICE_X5Y123_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D6 = CLBLM_R_X11Y128_SLICE_X15Y128_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A1 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A4 = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A6 = CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B1 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B4 = CLBLM_L_X10Y128_SLICE_X12Y128_DQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_DQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C3 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C4 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C5 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D4 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D5 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D6 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B6 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = CLBLM_R_X7Y124_SLICE_X8Y124_DQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = CLBLL_L_X4Y127_SLICE_X4Y127_DQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_A5Q;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AX = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = CLBLM_R_X7Y124_SLICE_X8Y124_DQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C5 = CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B4 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A2 = CLBLM_L_X10Y122_SLICE_X13Y122_B5Q;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D2 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D5 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D6 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = CLBLM_L_X8Y124_SLICE_X11Y124_CQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = CLBLM_L_X8Y122_SLICE_X11Y122_DQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_C5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = CLBLL_L_X4Y128_SLICE_X4Y128_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_AX = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = CLBLM_R_X13Y124_SLICE_X18Y124_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = CLBLL_L_X4Y127_SLICE_X5Y127_A5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = CLBLM_R_X5Y123_SLICE_X7Y123_A5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_A5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D5 = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A3 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A4 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A5 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B2 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B6 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C2 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C4 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C5 = CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D1 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D3 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D4 = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D6 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A1 = CLBLL_L_X4Y128_SLICE_X5Y128_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A3 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A5 = CLBLM_L_X12Y126_SLICE_X17Y126_DQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A6 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B1 = CLBLL_L_X4Y127_SLICE_X5Y127_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B2 = CLBLM_R_X7Y127_SLICE_X8Y127_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B3 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B5 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B6 = CLBLL_L_X4Y128_SLICE_X4Y128_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C1 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C2 = CLBLM_L_X8Y133_SLICE_X10Y133_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C6 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D2 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D3 = CLBLL_L_X4Y125_SLICE_X4Y125_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D4 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D5 = CLBLL_L_X4Y128_SLICE_X5Y128_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B3 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B4 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C5 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C6 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_CE = LIOB33_X0Y77_IOB_X0Y77_I;
endmodule
