module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y63_IOB_X0Y64_OPAD,
  output LIOB33_X0Y65_IOB_X0Y65_OPAD,
  output LIOB33_X0Y65_IOB_X0Y66_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AMUX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BQ;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CLK;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CMUX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A5Q;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C5Q;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CE;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CLK;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A5Q;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CLK;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B5Q;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C5Q;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D5Q;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CLK;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DQ;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CLK;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CLK;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D5Q;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DQ;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C5Q;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C5Q;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CE;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B5Q;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A5Q;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C5Q;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5Q;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D5Q;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CE;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A5Q;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B5Q;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C5Q;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CE;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D5Q;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CLK;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A5Q;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CLK;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A5Q;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AMUX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B5Q;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BMUX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BMUX;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CLK;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CLK;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B5Q;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BMUX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AMUX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CE;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CLK;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CE;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CLK;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CLK;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CMUX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DMUX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CE;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CLK;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CLK;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C5Q;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CE;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D5Q;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DMUX;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C5Q;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CMUX;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D5Q;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DMUX;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C5Q;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CMUX;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D5Q;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DMUX;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A5Q;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AMUX;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B5Q;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BMUX;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C5Q;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CMUX;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A5Q;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B5Q;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D5Q;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C5Q;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D5Q;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5Q;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5Q;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5Q;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5Q;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CE;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CE;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5Q;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5Q;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5Q;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5Q;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CE;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A5Q;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AMUX;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B5Q;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BMUX;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CMUX;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DMUX;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CE;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A5Q;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B5Q;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DMUX;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CE;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CE;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CLK;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A5Q;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CLK;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C5Q;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CLK;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CLK;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D5Q;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B5Q;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C5Q;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AMUX;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AX;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CE;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CLK;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CMUX;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CLK;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CLK;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AMUX;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BMUX;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AMUX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CE;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CLK;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CMUX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AMUX;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CMUX;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AMUX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BMUX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_CO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_CO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_DO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_DO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_DO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CLK;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CLK;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CLK;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B5Q;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C5Q;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CLK;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CLK;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_DO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AX;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_BO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CE;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CLK;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_DO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CLK;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CLK;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CLK;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CLK;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B5Q;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B5Q;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5Q;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5Q;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5Q;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5Q;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5Q;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5Q;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5Q;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CE;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5Q;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D5Q;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B5Q;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C5Q;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D5Q;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5Q;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_TQ;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y55_IOB_X0Y56_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.Q(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y123_SLICE_X1Y123_BO6),
.Q(CLBLL_L_X2Y123_SLICE_X1Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000080000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_CLUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_BQ),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00ee44aa00)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I4(LIOB33_X0Y53_IOB_X0Y54_I),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_CO6),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff00088008800)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AQ),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_AO5),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5fafaff5f5fafa)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_BLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_C5Q),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffaa00aa)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_ALUT (
.I0(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff780078ff780078)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_ALUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_BO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_CO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc000000cc000000)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50eeee4444)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_A5Q),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff600f688888888)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc5acc00)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_BO5),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.Q(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000300)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f00ff00c0c00000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_BLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.I4(LIOB33_X0Y57_IOB_X0Y58_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40aa000000ffff)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I4(LIOB33_X0Y57_IOB_X0Y58_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X4Y126_AO6),
.Q(CLBLL_L_X4Y126_SLICE_X5Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X5Y126_CO5),
.Q(CLBLL_L_X4Y126_SLICE_X5Y126_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X5Y126_AO6),
.Q(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X5Y126_BO6),
.Q(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.Q(CLBLL_L_X4Y126_SLICE_X5Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_DLUT (
.I0(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afafa0a0)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_CLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_C5Q),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_B5Q),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff010001ff300030)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffef00efffcf00cf)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_ALUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_BO5),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_BO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_CO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.Q(CLBLL_L_X4Y127_SLICE_X4Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afa0afa0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_DLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_C5Q),
.I1(LIOB33_X0Y63_IOB_X0Y63_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fafa0a0a)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006666ccccf0f0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_BQ),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a3a0a0a0a3a0)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_AO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y127_SLICE_X5Y127_DO6),
.Q(CLBLL_L_X4Y127_SLICE_X5Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaacfaaff)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_DLUT (
.I0(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I5(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aac0aaffaacc)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_DQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0f0f003000000)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I5(CLBLM_R_X5Y129_SLICE_X7Y129_A5Q),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00bb11aa00ea40)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_B5Q),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_CO5),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_BO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X4Y128_CO6),
.Q(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00a0a0f5f5)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_B5Q),
.I3(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000808ff000000)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_BLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_C5Q),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54aa00fe54)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_CO5),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_DO5),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_AO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_BO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_CO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_DO6),
.Q(CLBLL_L_X4Y128_SLICE_X5Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888dd88f5f5a0a0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_DQ),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_B5Q),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff55a0a0f5f5)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff6fffc0f060f0c)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_BLUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_DO6),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_A5Q),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdd00ddffd000d0)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_C5Q),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_CO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_DO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaff003a3a)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef000fe0efe0e)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_CLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_C5Q),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2c0e2f3e2)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I5(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaa0ccccfff0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_CO5),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_BO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_CO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff55ffffff)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_A5Q),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff990000ff99)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_BLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00eeeeff00ffff)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_ALUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_AO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_BO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_CO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_DO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cfacacacac)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y129_SLICE_X7Y129_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ff00cccc)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a8a8ff00fcfc)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_B5Q),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_BO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbfffbfafafffa)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_DO6),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_DO6),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccffaaccaacc)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_A5Q),
.I1(CLBLM_R_X3Y130_SLICE_X2Y130_A5Q),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fc54fc54)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_ALUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_D5Q),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_B5Q),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8000ffff0000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_CLUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff77ff80008000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_BLUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faaf0cc00ccff)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_DQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_BO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_CO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffc)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(CLBLM_R_X5Y133_SLICE_X6Y133_CQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_B5Q),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbebe1414ff55aa00)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_A5Q),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa00aacc)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_BLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_DQ),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00003c003c00)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_CO5),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_BO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_CO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_DO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffff3300)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_DLUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4b1e4fafa5050)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_C5Q),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaaf333)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_BLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa0caaf0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X6Y133_CQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_DQ),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_DLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_C5Q),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0aa00ee44)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I2(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_DQ),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa303c3c3c3c3c)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_BLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_C5Q),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ddf0dddddddddd)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_A5Q),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7f7fffffffff)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_BLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ff0000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_ALUT (
.I0(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_BO6),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_CO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a3b00330a0a0000)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00fc00fc)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_C5Q),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.I2(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcf00cfffc000c0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I5(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0fa50)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_ALUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_AO5),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300e2e2e2e2)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000fffc3330)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_DO6),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_BO6),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8d8d8dafaf0505)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a8a8ff00fcfc)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_BLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caac0aa0caac0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_DQ),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cccc0aa0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_DLUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AO6),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0c00000f0c0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_CO6),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeaafe54540054)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc5acc00ccf0cc00)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_B5Q),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_DQ),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800080008000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_DLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_AO6),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_CLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a000aa00aa00)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_BO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_CO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_DO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000bbb0bbb0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_DLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_DQ),
.I3(CLBLL_L_X4Y127_SLICE_X4Y127_D5Q),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0054545454)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_CLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_DQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfcf8fc0d0c080c)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ec20ff33fc30)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_C5Q),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_DO5),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_CO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_DO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd88dd8fafa5050)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_C5Q),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heefaeefa44504450)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa0faaccaa0c)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_B5Q),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb88888bb88bb8)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_C5Q),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_DO5),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_CO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_DO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaff00aaaa)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f055aaccccaaaa)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_DQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0acacafa0afa0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_BLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_DQ),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88b8b8b8b8)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_ALUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_CO5),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_DO5),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_CO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_DO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ffcc00cc)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_DLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_CO6),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88ddfafa5050)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_D5Q),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_C5Q),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300ffff3333)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_C5Q),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haacfaa03aafcaa30)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_B5Q),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_C5Q),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_BO5),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_CO5),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_CO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ffff6666ffff66)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_D5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30b8b8b8b8)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_CLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030de12de12)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_BLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_D5Q),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa33ff5a005a)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_BO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_CO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_DO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ffcc00ccff)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaffcc00ccff)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_CLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_C5Q),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc008bb88bb8)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_BLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50eeee4444)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_CO5),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_DO5),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_BO6),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_CO6),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_DO6),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bbbb88f3c0f3c0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_DLUT (
.I0(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ff3c003c)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaa330000aa33)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_CQ),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000a2a8a2a8)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I2(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_CO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_DO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaacccc)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_C5Q),
.I1(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_B5Q),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300e2e2e2e2)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_DQ),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22fcfc3030)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(RIOB33_X105Y123_IOB_X1Y124_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88bb88b888b8)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_CO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_DO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888e4e4e4e4)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cacacaca)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_C5Q),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e4e4ff00f0f0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.I2(CLBLM_L_X8Y129_SLICE_X11Y129_CQ),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf3aac0aaf3aac0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000000c)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_B5Q),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_DO6),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_B5Q),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_C5Q),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_DQ),
.I4(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_B5Q),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0a00000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfcfc0acacacac)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I1(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffee00005544)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfc0cfc0c)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I4(CLBLM_R_X7Y135_SLICE_X8Y135_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0ccaaccaacca0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_D5Q),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_D5Q),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_B5Q),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ccfffff0fc)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_CO6),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030ff30babaffba)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_DQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_DQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_B5Q),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_CO6),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00000ec20cc00)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_BLUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3131fffff5f5ffff)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I3(1'b1),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_CO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00cccc)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_B5Q),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11ee22f3c0f3c0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_CLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_D5Q),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0f505fa0a)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_BLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_D5Q),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y129_SLICE_X7Y129_C5Q),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaccaacc)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_ALUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_DQ),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_BO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_DO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaf05058d8d8d8d)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00eeeeff000e0e)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_C5Q),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ccccccf0f0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_B5Q),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0aa000000aa0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_DQ),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_BO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_CO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_DO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haafe0054aafe0054)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_DQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0a0f5e4f5e4)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_CQ),
.I2(CLBLM_L_X8Y135_SLICE_X11Y135_C5Q),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_D5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf303aaaafc0c)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cff0ff000f)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_CO5),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_DO5),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_BO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_CO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_DO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0acfc0cfc0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03fc30bbbb8888)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_B5Q),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf8fffc0a080f0c)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I5(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00d8d8ff00d8d8)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_BQ),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_CO5),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_BO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_CO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00e4e4e4e4)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_DQ),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_DQ),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0aaccf0ccf0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0c0c0cfc0c5c0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_BLUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf8fbf80b080b08)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_B5Q),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffffffffffff)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.I5(CLBLM_L_X8Y135_SLICE_X11Y135_BQ),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000044)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_CLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_AO6),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cfcfc0c0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050cc000000)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_CQ),
.I4(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_CO5),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_BO6),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_CO6),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_DLUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_BQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888ee44ee44)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafa3aca3ac)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefcee22223022)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff08ffff0000ffff)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffc000550015)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_ALUT (
.I0(CLBLM_L_X10Y126_SLICE_X12Y126_DQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_B5Q),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c000cc00cc00)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000e0eee0ee)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_CLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff6f0f60f060006)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_DO6),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DQ),
.I5(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacffcaaaa0330)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_ALUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_C5Q),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ee44fa50fa50)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecc3200fefe3232)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X10Y127_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008b00000088)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_DO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habaa0100aaaa0000)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_D5Q),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccff00cccc)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_CQ),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hce02ec20ec20ec20)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_ALUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AO6),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_AO5),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaaaa2a)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0fffff4f0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_D5Q),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_CQ),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccccaaccf0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_B5Q),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_B5Q),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_BO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_DO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00000aa00)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_DO6),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ffcc00ccff)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccf0ccf0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_BLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffde00deff120012)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_A5Q),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400f40004000400)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_CLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AO5),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_D5Q),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h08085d0800000000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_BLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_AO5),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_D5Q),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0503000305000000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_D5Q),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_DO5),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_DO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444f5a0f5a0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_D5Q),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4f5e4a0e4a0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00cacacaca)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_A5Q),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ec20ff33fc30)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_C5Q),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030ffff30303030)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaaabaaaaabbaaaa)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_CLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_AO6),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_B5Q),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3000ffff0022)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_BLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_C5Q),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_AO6),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaeaeffffffae)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_D5Q),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_CO6),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_DQ),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fffafffff5fffa)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_DLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_A5Q),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9000090000900009)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_CLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_C5Q),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeffeffffffff)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_DO6),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_DO6),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I5(CLBLM_L_X10Y128_SLICE_X12Y128_CO6),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_BO5),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5fafaff5f5fafa)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_B5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeffffffffe)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_BLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_DO6),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_DO6),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0fff000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_ALUT (
.I0(CLBLM_R_X7Y128_SLICE_X9Y128_D5Q),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_D5Q),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_BO5),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_BO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6f6f6ff6f6f6f6)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_DLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_DQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffafefffffaaee)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_CLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_DO6),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_CQ),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f033aa33aa33)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccaaccaa)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_B5Q),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_A5Q),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_CO5),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_BO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ffbaff3030baba)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_DLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_C5Q),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0f3eeee2222)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_CLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444ffaa5500)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeff2233ecfc2030)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_CO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808030008080300)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_C5Q),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.I3(CLBLM_R_X5Y129_SLICE_X7Y129_C5Q),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f033aa33aa33)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_C5Q),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.I2(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f00300cacacaca)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22fc30ee22ee22)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aaffff00aa00aa)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0fdfcf5f0fdfc)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_DO6),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_C5Q),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffaaafeee)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X13Y130_DO6),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_D5Q),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_CO6),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7ffffffff7)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_CO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff00aaaa)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I3(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf3fcf3fc)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fcfc)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f4b0f4b0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa000000880088)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_C5Q),
.I2(1'b1),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_D5Q),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a0affffcece)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_A5Q),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.I3(1'b1),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_CO6),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00bf00)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff2fffffff22)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_BO6),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_DQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fcfc3030)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_DQ),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaff88cc)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafff8fc0a0f080c)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_D5Q),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0ff00)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_C5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_CQ),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000f500a0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(1'b1),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaeefe00f0ccfc)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_DQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaa00320010)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_D5Q),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0cc000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_A5Q),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_D5Q),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_DO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e2e2e2e2)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_DQ),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54aa00fe54fe54)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfeece33032202)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_BLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04ea40ea40ea40)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_DO5),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_CO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_DQ),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_AQ),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0c0aaaaffcc)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_CLUT (
.I0(CLBLM_L_X8Y129_SLICE_X11Y129_D5Q),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_CQ),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaff88cc)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff505fa0af000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_CQ),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_BO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffefee)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_DLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_C5Q),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_D5Q),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cccccc00cc6ccc)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_B5Q),
.I2(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaa5000feee5444)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_BO6),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdc1310cfcc0300)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_ALUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_BO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_DO5),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ffffffffffffff)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_B5Q),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_B5Q),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I5(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fef001000300030)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_BLUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_DO6),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffff5a005a)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_ALUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.I1(1'b1),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_B5Q),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_BO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_CO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f7ffffffffffff)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_DLUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CQ),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a0aca0aca0ac)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_CLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000beee1444)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_B5Q),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffcc5accf0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_ALUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_CO6),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffffff0c0c0c0c)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_DLUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa003cc0c0c0c0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_CLUT (
.I0(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_A5Q),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f055dd)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_C5Q),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f8f80808)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_ALUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_D5Q),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_AO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_BO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff7fffffff)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_DLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4a00f0f0f0f)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc30aaaacc00)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_BLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_C5Q),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.I3(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfe3032ccce0002)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_ALUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.I4(CLBLM_L_X8Y135_SLICE_X11Y135_BQ),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_CO6),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.Q(CLBLM_L_X10Y136_SLICE_X13Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.Q(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.Q(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffffffffff)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_DLUT (
.I0(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0400040a0a0a0a)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c0c0ff00e2e2)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_BLUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AO6),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000505ff003535)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_ALUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_DO6),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h007f7f7f00ffffff)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_BLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32fe32ce02ce02)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_ALUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_CO6),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_AO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_BO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_CO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc3333cccc3333)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc3cccca5a6a5a5)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_BLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_B5Q),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_BQ),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_DO6),
.I3(CLBLM_L_X12Y124_SLICE_X16Y124_CQ),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00110000f0ff0f00)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_ALUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_B5Q),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_BQ),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_DO6),
.I3(CLBLM_L_X12Y124_SLICE_X16Y124_CQ),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffdff)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_CLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffffffbffff)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111005000000050)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_DLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffeffffff)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_BLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3fcaaaa0000)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafefafefafeffff)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_DLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_CO6),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_DQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_AO6),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbffff)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffff)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7fffffdff)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_BO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_CO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'habaaafafabaaabaa)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_DLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdf8f80d0d0808)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_CLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0cccc)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccc0fff0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_ALUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000020f)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_AO6),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_BO6),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_DO6),
.I5(CLBLM_R_X11Y130_SLICE_X15Y130_BO6),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeffffffff77)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffffffefffff)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffbfffff)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_ALUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_AO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfefffffccee)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_DLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_DO6),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_DO6),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008b00000088)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_CLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55a8b8b8b8b)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_BLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa00ccccfafa)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010111110100000)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_DLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddfddcccccfcc)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_CLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_AO6),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_CO6),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff00ac)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_AO6),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff0cffffffae)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_ALUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_BO6),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X16Y129_AO6),
.Q(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.Q(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfff0fffccff00)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_CO6),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I5(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200030002000000)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_C5Q),
.I1(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff0c00fc000c)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecc3200fefe3232)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfefecccceeee)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I2(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_AO5),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeefffffffe)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_CLUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_AO6),
.I1(CLBLM_L_X12Y128_SLICE_X17Y128_DO6),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_DO6),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050405)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_BLUT (
.I0(CLBLM_R_X11Y129_SLICE_X15Y129_DO6),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_CO6),
.I2(CLBLM_R_X11Y129_SLICE_X15Y129_BO6),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_CO6),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_CO6),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0cff0caeaeffae)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X17Y130_DO6),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_CQ),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_AO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_BO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00aaaaff00)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044004500440044)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_CLUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_DO6),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_AO5),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_DO6),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_BO6),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffaa00aa)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aaf0aaf0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010000055100000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_DLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_D5Q),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000a0a00cc0ace)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I2(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff0cffffffae)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_D5Q),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_CO6),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_AO6),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_AO6),
.I5(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffffb)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_ALUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_CQ),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699696696996)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_DLUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_BO6),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff01310000)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_AO5),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_DO6),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff04ff40ff44)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_BLUT (
.I0(CLBLM_L_X12Y133_SLICE_X17Y133_DO6),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_BO6),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_ALUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_D5Q),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_BO6),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I4(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I5(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y131_SLICE_X18Y131_BO5),
.Q(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f4b5a000f445a)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_DLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I1(CLBLM_R_X13Y131_SLICE_X18Y131_DO6),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_DO6),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_DO6),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_CO6),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0022222f22)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffaa)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_BLUT (
.I0(CLBLM_L_X12Y129_SLICE_X16Y129_DO6),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.I3(CLBLM_L_X12Y130_SLICE_X17Y130_BO6),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_BO6),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccdccccdcddcccc)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_ALUT (
.I0(CLBLM_L_X12Y133_SLICE_X17Y133_CO6),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I4(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_DO5),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_CO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_DO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaff0ff000)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X18Y130_AO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_CQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f5f5c4c4)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_CLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_B5Q),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heedd2211dedd1211)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_BLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_L_X8Y128_SLICE_X10Y128_D5Q),
.I4(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaaf0fc)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_ALUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y132_SLICE_X15Y132_A5Q),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5055505510111011)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_DLUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_R_X13Y133_SLICE_X18Y133_AO6),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaaaaaa)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_DO6),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_BO6),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc040cc44f050ff55)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_BLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_DQ),
.I1(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_AO6),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I5(RIOB33_X105Y143_IOB_X1Y143_I),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff22ff2222)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_ALUT (
.I0(LIOB33_X0Y51_IOB_X0Y52_I),
.I1(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I3(CLBLM_R_X13Y133_SLICE_X18Y133_BO6),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_CO5),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_AO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_BO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_CO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbfffffff0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_DLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0f5f50505)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_CLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.I4(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccffcccc)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff320032ff300030)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.Q(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.Q(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f0f0fff5fff0)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_DLUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.I1(1'b1),
.I2(CLBLM_L_X12Y134_SLICE_X17Y134_CO6),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(CLBLM_R_X13Y133_SLICE_X18Y133_AO6),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff55dd00cc)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_CLUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.I1(RIOB33_X105Y139_IOB_X1Y140_I),
.I2(1'b1),
.I3(CLBLM_R_X13Y133_SLICE_X18Y133_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(CLBLM_L_X12Y133_SLICE_X17Y133_BO6),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000044440f004f44)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I1(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0ddd0dd0000d0dd)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_ALUT (
.I0(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I1(CLBLM_R_X13Y133_SLICE_X18Y133_AO6),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_AO6),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.Q(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbbbb8b8b8)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X13Y134_SLICE_X18Y134_BO6),
.I3(RIOB33_X105Y139_IOB_X1Y139_I),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_DO6),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaaaaaf0f00000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y139_IOB_X1Y140_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y141_I),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000222233000000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I1(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I2(1'b1),
.I3(RIOB33_X105Y139_IOB_X1Y139_I),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff888f888f888)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_BLUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_BQ),
.I2(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(RIOB33_X105Y143_IOB_X1Y144_I),
.I5(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05040100fbfbfbfb)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I3(RIOB33_X105Y143_IOB_X1Y144_I),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_BO6),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa00aa00aa)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.I3(CLBLL_L_X2Y123_SLICE_X1Y123_BQ),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_AQ),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa30c030c0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.I2(LIOB33_X0Y53_IOB_X0Y54_I),
.I3(CLBLL_L_X2Y123_SLICE_X1Y123_CO5),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff007d7d7d7d)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff30ff3000300030)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_BQ),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066006600)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000078ff78ff)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_AQ),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_D5Q),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000005)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_ALUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_BO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_C5Q),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I5(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.Q(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f000000fffb)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_CLUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_C5Q),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_D5Q),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000c000f0000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_BLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_A5Q),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffff0033)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_ALUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_BO5),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_CO5),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_BO6),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.Q(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y122_I),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0fff000)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfcecfc31302030)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_AQ),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_CQ),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_BQ),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X3Y127_AO5),
.Q(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.Q(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.Q(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffefefffff)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_DLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_C5Q),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000b0b00000b0a)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_CLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I2(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_C5Q),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30ff33fc30fd31)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_BLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_D5Q),
.I5(CLBLM_R_X3Y127_SLICE_X3Y127_CO6),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaf0f0cccc)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_D5Q),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_D5Q),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_DO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_CO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_BO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_AO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.Q(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_DO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_CO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000cc00440044)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_BLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_C5Q),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_BQ),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_BO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff00ff30ff00)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_ALUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_C5Q),
.I3(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_BQ),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_AO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.Q(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X2Y129_BO6),
.Q(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fff7f00800000)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f8f2f802080208)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I1(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y130_SLICE_X2Y130_BO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_B5Q),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heecc2200ceec0220)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_C5Q),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_AO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_BO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_CO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.Q(CLBLM_R_X3Y129_SLICE_X3Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fccf0cc0fccf0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(LIOB33_X0Y59_IOB_X0Y60_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdd00ddff000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_CQ),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000dd0000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_BLUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_CO6),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_BQ),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00bbbbb0b0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_BQ),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.Q(CLBLM_R_X3Y130_SLICE_X2Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X2Y130_AO6),
.Q(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee444430003000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000082828282)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.Q(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32fe32dc10dc10)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_ALUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_D5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050505050505050)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y127_SLICE_X2Y127_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_AO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf5fa0a05f5fa0a0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_CLUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I1(LIOB33_X0Y55_IOB_X0Y55_I),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_A5Q),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccaaaaf333)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I2(LIOB33_X0Y55_IOB_X0Y55_I),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aaf0aaf0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.I2(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdefc123000ff00ff)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_ALUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(LIOB33_X0Y59_IOB_X0Y60_I),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_BO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_CO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_DO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff1c001c)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ddddff00d0d0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_CLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_B5Q),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff0055dddd8888)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff007070f0f0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_ALUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_DQ),
.I1(LIOB33_X0Y59_IOB_X0Y60_I),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_BO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff000000ff00)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafacff0ff000)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_C5Q),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000404ff004040)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_CO6),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7bff7bffdeffde)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_DLUT (
.I0(CLBLL_L_X4Y124_SLICE_X5Y124_A5Q),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_DQ),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.I3(CLBLL_L_X4Y124_SLICE_X5Y124_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y127_SLICE_X2Y127_BQ),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff6ffffffff6)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_D5Q),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_CO6),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.I5(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acacacaca)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_BLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I1(CLBLL_L_X4Y124_SLICE_X5Y124_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0f0cccc)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h880088005fffffff)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_CO6),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbaaee00110044)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I5(CLBLL_L_X4Y127_SLICE_X5Y127_AQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a3a3a3a0a0a0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_B5Q),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_CO6),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a8a8ff00fcfc)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_CO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000100010001)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_DLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_C5Q),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_DO6),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y61_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5a0f5a0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fa0afa0a)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_BLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_DQ),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00de12cc00de12)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_CO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_DO6),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I5(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0eeee4444)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ff606fc0c)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fafaff003232)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_B5Q),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8822882244114411)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_D5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5ff5f5afaffafa)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_D5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff5ff5)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14be14ffaa5500)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_CO6),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_DO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaf0505dddd8888)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0ac0c0cfc0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_C5Q),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_A5Q),
.I4(CLBLM_L_X8Y134_SLICE_X11Y134_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0cc0000f0cc)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aa33aa30)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I1(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_DO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f3f3fcfc)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_BO6),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30eeee2222)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(RIOB33_X105Y123_IOB_X1Y123_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_DQ),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a3aca0a0acac)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_CQ),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_BO6),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdefccccc12300000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_C5Q),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_CO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaf0f0cccc)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afff00f00)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_CLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_A5Q),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_D5Q),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfef55551545)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AO6),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88d8d8dd88dd88)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_CO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_DO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc55f055f055)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_DLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc55ff550055)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aacc55ccaa)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_BLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_C5Q),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0ffaa5500)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_CO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_DO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfc3130ecfc2030)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_C5Q),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8bb8b888888)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000000f000f)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_CO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330033aa33aa33)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafa0f0f0a0a)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_BO6),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cfafa0afa0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7fffffffff)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc6ccccccccc)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00fff000f0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_CQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5a0dd88dd88)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_CO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_C5Q),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_DQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaaaaa3c3c)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aabf0015)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I4(CLBLM_L_X8Y134_SLICE_X10Y134_D5Q),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffe0f0e0f0e)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y127_SLICE_X2Y127_B5Q),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_AO5),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_DO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222e2e2e2e2)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0ac5cac5ca)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_C5Q),
.I4(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff6fff60f060f06)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_BLUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_DO6),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfafa0a0a)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_DO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_D5Q),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_AO5),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_CO5),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa0fccf0ccf0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_DLUT (
.I0(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaff660066)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_CLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dddd88e4e4e4e4)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ffaa5500)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_DO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ccaaf0aaf0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0fa50fa50)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_DQ),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_A5Q),
.I4(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddd8d88d88888)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I5(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888ddd8ddd8)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_DQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0bbbb8888)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404f303f404)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_CLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_B5Q),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_AO6),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcf0fc0f0c000c)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff338888bbbb)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_AO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_BO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_CO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_DO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccc44ee)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_DLUT (
.I0(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff660066f0fff000)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00afaf8c8c)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_BLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_D5Q),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_A5Q),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888b8b8b8bbb8b8)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_ALUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I5(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_AO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0cc00ee22)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_CLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_D5Q),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eebbf0f0eeee)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_CO6),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff400f4ffb000b0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555beee1444)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_B5Q),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ce02ee22fe32)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_ALUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_CQ),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a0a0a0a0a)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_D5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00000000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_B5Q),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_C5Q),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaf0ccf0cc)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_ALUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_C5Q),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_AO5),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_BO5),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaaaaa0f0f)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_DQ),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaaaaaf0f0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800095559555)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_CLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f0040000550055)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_BLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b888b88b888b888)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333388d8d888)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I2(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I3(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00000000000)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff20200000)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f03300f0f0bbaa)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_BLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_DQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_CO6),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffcccc5a5a)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_ALUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_DO6),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff00ff)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f8f8f8f8f800)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_DO6),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0aca3a0a0a0a0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f10301f3f00300)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_DO6),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_AO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_DLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_CLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf033aaaaf0cc)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_A5Q),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_B5Q),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4a0f5f5a0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_C5Q),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000000000)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I4(1'b1),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaffffffff55aa)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_D5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafff0aaaa3330)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I1(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5b1e4e4e4)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_B5Q),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_DO6),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff003030)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff03aaaaff03)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_B5Q),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_DO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_C5Q),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ff55ee44aa00)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030de12de12)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0faccccf050)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_C5Q),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca0f5f5f5)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0ccfc0cfc0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabbee00001144)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_BO6),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I5(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44af05fa50)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_DO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0a0afa0af)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_DLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333aaaaf0f0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_DQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habae0104abae0104)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_B5Q),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_DO6),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_D5Q),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdceffcccccccccc)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_DO6),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I5(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_CLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0000005ff5affa)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_C5Q),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_DQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000003fffffff)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_DO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafffafaa05550500)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_B5Q),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dd118888bbbb)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_D5Q),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff6c0000006c)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y127_SLICE_X3Y127_AQ),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_CQ),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa30aa30)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_DO5),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_BO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_CO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_DO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00fff0f01111)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_DLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(CLBLL_L_X4Y127_SLICE_X5Y127_DQ),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f50505cfcfc0c0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_CLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eefff0f04400)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hde12de12ffcc3300)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_CO5),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_DO5),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_CO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee448888dddd)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fa050acacacaca)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_C5Q),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000cacacaca)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I4(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e4e4ff00f0f0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_C5Q),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habaaabaa01000100)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.I3(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfff00c0c0f00)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044faee5044)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_AQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_CO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_DO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888ddddd8d8)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacafa0afa0a)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50e4e4e4e4)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_B5Q),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddddd888888888)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_BQ),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_C5Q),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff7fffff)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffe3f3fffff)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_BQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffa0f0a0f0a)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_CO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_DO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff00aaaa)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_DLUT (
.I0(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_CLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_CQ),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500b1e4b1e4)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_C5Q),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_BQ),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000048c048c0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_DO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500f5a0f5a0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_A5Q),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haffa0550d8d8d8d8)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_A5Q),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_B5Q),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0c5c5)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0cc0aaaa0cc0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeeffffffee)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_C5Q),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbebe1414dd88dd88)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00acacacac)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaa0ccccfff0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_DQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_BO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_CO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff55ff55ff)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f0ccaaf0aaf0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X2Y130_AQ),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff202f202f202)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_B5Q),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_AO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888bbb8bbb8)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_D5Q),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_DQ),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_DQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbffbbcfcfc0c0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0fff000f0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fa0afa0a)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_BO5),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_CO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_DO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccfaccaf)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_D5Q),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff2300000023)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_D5Q),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccf0ccf0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_BLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_B5Q),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_CO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa03303030)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_B5Q),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_CO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11ee44e4e4e4e4)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_BQ),
.I4(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fafa5050)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00fff300f3)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0fcc00ccf0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_BO5),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_CO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc0ccc0c)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcfcacfca)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_CLUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_DQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacafff00f00)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb88bb88bb)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_ALUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_DO5),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_CO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afa0afa0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_DLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000abaf0105)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff558888dddd)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5555ff00aaaa)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_AO6),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_BO6),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_CO6),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_DO6),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccaaccaa)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff0fff0f)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_CLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3fc0000f3fc)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0acca0cca0cca0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_DQ),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_AO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_AO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_BO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00c033333333)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_B5Q),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff606ff0ffc0c)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_CLUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444faee5044)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_DQ),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_D5Q),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeff4455eafa4050)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_A5Q),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_BO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_DLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ef00df30303030)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_CLUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_C5Q),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a3acafafa3ac)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_BLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_CO5),
.I5(CLBLM_L_X10Y125_SLICE_X13Y125_A5Q),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5a005aff000000)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I5(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_BO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h880000003fffffff)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff006c6c0000)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_CLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_DQ),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff606000006060)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I2(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f80208faf00a00)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e0000000e0000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_ALUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_AO6),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccccffffcccc)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_DO5),
.I2(1'b1),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_BO5),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ff55aa00)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_C5Q),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I4(CLBLL_L_X4Y130_SLICE_X4Y130_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaf0f0cccc)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_BO5),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f00000)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050dd88dd88)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0f6f60f000606)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_ALUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_B5Q),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AO5),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_BO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_CO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ffaa00aa)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_CLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888cfcc0300)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X4Y127_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ffaa00aa)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0aff3bff0aff0a)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_DLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_CO6),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010b0100000a000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AO5),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_DQ),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3030ffff3075)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_BLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_A5Q),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_AO6),
.I5(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200000022a000a0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_A5Q),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0fcfffff00cc)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_B5Q),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_DO6),
.I5(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h505050dc50505050)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_CLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_CQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_DQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h220020205555ffff)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_C5Q),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_BO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0203020000000000)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_DLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_B5Q),
.I1(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_BQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffaaaeaeffae)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_CLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_CO6),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_C5Q),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I3(CLBLM_R_X5Y129_SLICE_X7Y129_A5Q),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00dddd8888)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3330aaaa3330)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_ALUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_B5Q),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_AO5),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfbaafabbfbaafa)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_DLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a020a0208000800)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_CLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_A5Q),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a4e000000440000)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_BLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_D5Q),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0ccf0cc)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f2f2fff0fff2)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_C5Q),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_BO6),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_B5Q),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0aceceff0affce)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_AO6),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_AO5),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2fff2f2f22ff2222)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_B5Q),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AO6),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_AO5),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I5(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32ff33dc10cc00)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_CQ),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_BO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5ff5f5afaffafa)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_DQ),
.I5(CLBLM_R_X5Y129_SLICE_X7Y129_A5Q),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0fff000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_DQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaffaa00aa)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccfff000f0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_C5Q),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeffeeeeeeee)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_DLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f5f3f0f77553300)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_CLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_C5Q),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001500000005)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_DO6),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_DO6),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_CO6),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_DO6),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_DO6),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3bff0a3b3b0a0a)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_ALUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_B5Q),
.I1(CLBLM_L_X12Y127_SLICE_X17Y127_AO6),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.I3(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00cfcc0f00cfcc)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I2(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_BQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaeaeffff0c0c)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_CLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_C5Q),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_DO6),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffa)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_BLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_DO6),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_CO6),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffc000000fc)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff33bbffff00aa)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_CO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_DO6),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22f2ffff22f222f2)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_CLUT (
.I0(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.I2(CLBLM_L_X8Y128_SLICE_X11Y128_C5Q),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h44f444f4ffff44f4)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_BLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_CO6),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_A5Q),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_A5Q),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffccfffdffcc)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_CO6),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_BO6),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_BO6),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030ff303030ff30)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_CQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff22f2)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_CLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I1(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_BO6),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I2(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf222f222fffff222)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_BQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X15Y130_AO5),
.Q(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X15Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fa005000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_DLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I4(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000030200000002)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_CLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I1(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffeeffefefeeee)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.I3(CLBLM_L_X12Y130_SLICE_X17Y130_AO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_CQ),
.I5(CLBLM_R_X11Y130_SLICE_X15Y130_A5Q),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff003388bb88bb)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5ccf5cca0cca0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd800d8ffd800d8)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_CQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef40e04fef40e04)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888ddd8ddd8)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_D5Q),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I5(CLBLL_L_X4Y127_SLICE_X4Y127_CQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_BQ),
.Q(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.Q(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcffdcdcdcffdc)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.I1(CLBLM_R_X11Y130_SLICE_X15Y130_DO6),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_DQ),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffbfff)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbffffffff7ffff)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdffffffffe)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X14Y132_AO6),
.Q(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffee)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_DLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ffbbff00ffaa)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.I5(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff5dff0c)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaa0ff0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_DQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.Q(CLBLM_R_X11Y132_SLICE_X15Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X15Y132_BO5),
.Q(CLBLM_R_X11Y132_SLICE_X15Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X15Y132_AO6),
.Q(CLBLM_R_X11Y132_SLICE_X15Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.Q(CLBLM_R_X11Y132_SLICE_X15Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cc4400008800)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_DLUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I2(1'b1),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_D5Q),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfffffcfc)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_BO6),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_AO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_CO6),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888a0f5a0f5)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_CQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0f5aaff0055)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_C5Q),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_DQ),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_DO5),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_DO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaf0ccf0cc)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_DLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc00aaaafcfc)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_CQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc540000fc54)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_C5Q),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_DO5),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_AO6),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_BO6),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_CO6),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_DO6),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0f0ccf0cc)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbe00beff140014)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_CLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_C5Q),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_B5Q),
.I5(CLBLM_R_X11Y133_SLICE_X15Y133_D5Q),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f1fcfc04010c0c)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_BLUT (
.I0(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffa500000fa50)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_ALUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_CO5),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_BO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_CO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0d2f033003300)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_DLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500dd88dd88)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacafff00f00)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_BO6),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaefaaa54045000)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_CO6),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_BO6),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_A5Q),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.Q(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f099cc)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_C5Q),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff000c0c)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_CO6),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_BO6),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.Q(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_B5Q),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I2(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_B5Q),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00007fff0000ffff)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_B5Q),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f5f5f5f00ffffff)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_ALUT (
.I0(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.Q(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccf0ccf0)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y137_SLICE_X14Y137_AO6),
.Q(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0203ffff0303ffff)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_DQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_B5Q),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_CLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002000000)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5155555555555555)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_ALUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005500ff00ff00)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_B5Q),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa33c0c0c0c0)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_A5Q),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbffffffff)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_DLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbffff)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_CLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001030000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccff51004000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_CLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I5(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3fffffffffffff)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffffffffff)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I2(CLBLL_L_X4Y128_SLICE_X5Y128_C5Q),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_CQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_B5Q),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcefffdcc)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_CO6),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_DO6),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_DO6),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h111f1111000f0000)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_CLUT (
.I0(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.I4(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I5(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff7350)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_AO6),
.I5(CLBLM_R_X11Y129_SLICE_X14Y129_CO6),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500f5f0ddccfdfc)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_C5Q),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0f0fffff)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_BLUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f2f3f2f3)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_DLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I1(CLBLM_L_X12Y130_SLICE_X17Y130_CO6),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccfcccccccfcf)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I4(CLBLM_R_X13Y134_SLICE_X18Y134_AO5),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h11001f0f11001100)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_BLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.I1(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I3(LIOB33_X0Y51_IOB_X0Y51_I),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff700000400)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_CO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_AO5),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff20ff2a)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_CLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I1(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I5(CLBLM_R_X11Y125_SLICE_X15Y125_BO6),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699669696996)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_DO6),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_BO6),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I5(CLBLM_R_X13Y130_SLICE_X18Y130_CO6),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeeefffffefe)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_BO6),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_BO6),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I5(CLBLM_R_X13Y131_SLICE_X18Y131_CO6),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccecfcecf)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_CLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_CO6),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_BO6),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500373305000500)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_BLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.I1(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I5(RIOB33_X105Y141_IOB_X1Y141_I),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbddfbf8f8d8f8)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I4(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cf00cc00dd00cc)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_DLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.I4(CLBLM_R_X13Y132_SLICE_X19Y132_CO6),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_DO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccceccdfcc)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_CLUT (
.I0(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_DO6),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AQ),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_CO6),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffffc0c0cfcf)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_B5Q),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_BO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7ffffefff)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_DO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fffafff0f0fafa)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(1'b1),
.I2(CLBLM_R_X13Y133_SLICE_X18Y133_BO5),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I4(CLBLM_R_X13Y133_SLICE_X18Y133_BO6),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_CO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1511050011110000)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I1(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_BO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaeabafa)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.I2(CLBLM_R_X13Y132_SLICE_X19Y132_DO6),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I5(CLBLM_R_X13Y131_SLICE_X19Y131_CO6),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f0a0f0aaffaaff)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_DLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I1(1'b1),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.I3(RIOB33_X105Y145_IOB_X1Y145_I),
.I4(1'b1),
.I5(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hceffcececeffcece)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_CLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I1(CLBLM_R_X13Y133_SLICE_X18Y133_AO5),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I3(CLBLM_R_X13Y133_SLICE_X18Y133_BO6),
.I4(RIOB33_X105Y137_IOB_X1Y138_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h003000ba000000aa)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y138_I),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.I4(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040004400500055)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_ALUT (
.I0(CLBLM_R_X13Y133_SLICE_X18Y133_AO5),
.I1(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.I2(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y145_I),
.I5(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb0000bbbbbbbb)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_DLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000b0000000b000b)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_CLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X13Y133_SLICE_X18Y133_BO5),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_BO6),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3bbbbbbbb)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_DO6),
.I1(CLBLM_R_X11Y132_SLICE_X15Y132_B5Q),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f1f155ff55ff)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_ALUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_B5Q),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0f0f0f0f)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y132_SLICE_X15Y132_CO6),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_DO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaaf000f000)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_CLUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_CO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcffff0c000808)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_BLUT (
.I0(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_BO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f7f7f70c080400)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I2(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I3(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_AO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_DO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcf0f0fffff)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_CO6),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_B5Q),
.I3(1'b1),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_BO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55f5f5f5f5)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_ALUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_AO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ff00f0f00000)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y145_I),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I5(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_DO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ffa0a0a0a0a0)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(1'b1),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_CO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffee)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_BLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.I1(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_R_X13Y133_SLICE_X18Y133_CO6),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff000c000a0)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_D5Q),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_AO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_DO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_CO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_BO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_AO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y125_IOB_X1Y125_I),
.I2(1'b1),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(1'b1),
.I5(RIOB33_X105Y127_IOB_X1Y127_I),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y64_OBUF (
.I(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.O(LIOB33_X0Y63_IOB_X0Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y65_OBUF (
.I(CLBLM_R_X7Y123_SLICE_X8Y123_DO6),
.O(LIOB33_X0Y65_IOB_X0Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y66_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.O(LIOB33_X0Y65_IOB_X0Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X4Y125_SLICE_X5Y125_CQ),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X4Y126_SLICE_X5Y126_CQ),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X4Y130_SLICE_X4Y130_D5Q),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLM_R_X7Y126_SLICE_X8Y126_DQ),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X4Y126_SLICE_X5Y126_C5Q),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X7Y128_SLICE_X9Y128_DQ),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLM_R_X3Y127_SLICE_X3Y127_A5Q),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_R_X5Y127_SLICE_X6Y127_D5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X7Y132_SLICE_X8Y132_A5Q),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X9Y131_C5Q),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X11Y124_SLICE_X15Y124_B5Q),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_L_X10Y125_SLICE_X13Y125_A5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X7Y127_SLICE_X9Y127_DQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y131_SLICE_X11Y131_B5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X11Y133_SLICE_X14Y133_D5Q),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y75_SLICE_X0Y75_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X5Y127_BQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_L_X8Y134_SLICE_X11Y134_C5Q),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X6Y133_C5Q),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X4Y131_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X2Y131_AO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(CLBLM_R_X5Y129_SLICE_X6Y129_D5Q),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(CLBLL_L_X4Y127_SLICE_X4Y127_AQ),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(CLBLM_R_X5Y136_SLICE_X7Y136_AO6),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(CLBLM_R_X7Y135_SLICE_X9Y135_DO5),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(CLBLM_L_X8Y135_SLICE_X10Y135_BO6),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(CLBLM_R_X7Y132_SLICE_X8Y132_DO6),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(1'b1),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X5Y131_C5Q),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(1'b1),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X8Y132_SLICE_X11Y132_C5Q),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X8Y131_SLICE_X11Y131_D5Q),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X3Y128_SLICE_X3Y128_AQ),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X5Y136_SLICE_X7Y136_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X4Y131_CO6),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X3Y131_A5Q),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_R_X7Y132_SLICE_X8Y132_DO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_R_X11Y136_SLICE_X14Y136_DO6),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X8Y136_SLICE_X10Y136_BO6),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y133_SLICE_X19Y133_BO5),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X13Y133_SLICE_X18Y133_DO6),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y133_SLICE_X19Y133_AO6),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X13Y132_SLICE_X19Y132_BO6),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X13Y133_SLICE_X19Y133_AO5),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X13Y131_SLICE_X18Y131_BO6),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_R_X13Y132_SLICE_X19Y132_AO5),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X13Y133_SLICE_X19Y133_BO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(1'b1),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B = CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C = CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D = CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A = CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B = CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C = CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D = CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_AMUX = CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_CMUX = CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A = CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B = CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_AMUX = CLBLL_L_X4Y124_SLICE_X5Y124_A5Q;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A = CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A = CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_AMUX = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_BMUX = CLBLL_L_X4Y125_SLICE_X5Y125_BO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_CMUX = CLBLL_L_X4Y125_SLICE_X5Y125_C5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_AMUX = CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_BMUX = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_AMUX = CLBLL_L_X4Y126_SLICE_X5Y126_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_CMUX = CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A = CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B = CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_BMUX = CLBLL_L_X4Y127_SLICE_X4Y127_B5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_CMUX = CLBLL_L_X4Y127_SLICE_X4Y127_C5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_DMUX = CLBLL_L_X4Y127_SLICE_X4Y127_D5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A = CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B = CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C = CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D = CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_CMUX = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A = CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B = CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_CMUX = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_DMUX = CLBLL_L_X4Y128_SLICE_X5Y128_D5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A = CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_CMUX = CLBLL_L_X4Y129_SLICE_X5Y129_C5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_DMUX = CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_CMUX = CLBLL_L_X4Y130_SLICE_X4Y130_C5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_DMUX = CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_BMUX = CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_AMUX = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_BMUX = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_CMUX = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B = CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_CMUX = CLBLL_L_X4Y132_SLICE_X4Y132_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_AMUX = CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_BMUX = CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CMUX = CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A = CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B = CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A = CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_AMUX = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A = CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CMUX = CLBLM_L_X8Y125_SLICE_X10Y125_C5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A = CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_AMUX = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_DMUX = CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_AMUX = CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_BMUX = CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A = CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A = CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B = CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_DMUX = CLBLM_L_X8Y127_SLICE_X10Y127_D5Q;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A = CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B = CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_CMUX = CLBLM_L_X8Y127_SLICE_X11Y127_C5Q;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_DMUX = CLBLM_L_X8Y127_SLICE_X11Y127_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A = CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B = CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C = CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_CMUX = CLBLM_L_X8Y128_SLICE_X10Y128_C5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_DMUX = CLBLM_L_X8Y128_SLICE_X10Y128_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A = CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B = CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_AMUX = CLBLM_L_X8Y128_SLICE_X11Y128_A5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_BMUX = CLBLM_L_X8Y128_SLICE_X11Y128_B5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_CMUX = CLBLM_L_X8Y128_SLICE_X11Y128_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_AMUX = CLBLM_L_X8Y129_SLICE_X10Y129_A5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_BMUX = CLBLM_L_X8Y129_SLICE_X10Y129_B5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CMUX = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_DMUX = CLBLM_L_X8Y129_SLICE_X10Y129_D5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_CMUX = CLBLM_L_X8Y129_SLICE_X11Y129_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_DMUX = CLBLM_L_X8Y129_SLICE_X11Y129_D5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_BMUX = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CMUX = CLBLM_L_X8Y130_SLICE_X10Y130_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_DMUX = CLBLM_L_X8Y130_SLICE_X10Y130_D5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_CMUX = CLBLM_L_X8Y130_SLICE_X11Y130_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_DMUX = CLBLM_L_X8Y130_SLICE_X11Y130_D5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_AMUX = CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_BMUX = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_DMUX = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_AMUX = CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_BMUX = CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_AMUX = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_BMUX = CLBLM_L_X8Y132_SLICE_X11Y132_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CMUX = CLBLM_L_X8Y132_SLICE_X11Y132_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_BMUX = CLBLM_L_X8Y133_SLICE_X10Y133_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_DMUX = CLBLM_L_X8Y133_SLICE_X10Y133_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_AMUX = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A = CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_AMUX = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_CMUX = CLBLM_L_X8Y134_SLICE_X10Y134_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_DMUX = CLBLM_L_X8Y134_SLICE_X10Y134_D5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_CMUX = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_DMUX = CLBLM_L_X8Y134_SLICE_X11Y134_D5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A = CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_AMUX = CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_BMUX = CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_CMUX = CLBLM_L_X8Y135_SLICE_X11Y135_C5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_DMUX = CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_AMUX = CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A = CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B = CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_DMUX = CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_BMUX = CLBLM_L_X10Y125_SLICE_X12Y125_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A = CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_AMUX = CLBLM_L_X10Y125_SLICE_X13Y125_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_BMUX = CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A = CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CMUX = CLBLM_L_X10Y126_SLICE_X12Y126_C5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A = CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B = CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C = CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_BMUX = CLBLM_L_X10Y127_SLICE_X12Y127_B5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_DMUX = CLBLM_L_X10Y127_SLICE_X12Y127_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A = CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_DMUX = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_AMUX = CLBLM_L_X10Y128_SLICE_X13Y128_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_DMUX = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B = CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_AMUX = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_BMUX = CLBLM_L_X10Y129_SLICE_X12Y129_B5Q;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A = CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_CMUX = CLBLM_L_X10Y129_SLICE_X13Y129_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_BMUX = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CMUX = CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_AMUX = CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_DMUX = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_AMUX = CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_BMUX = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CMUX = CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A = CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A = CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_DMUX = CLBLM_L_X10Y133_SLICE_X13Y133_D5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A = CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B = CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A = CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_BMUX = CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_AMUX = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_CMUX = CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_DMUX = CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_AMUX = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CMUX = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_DMUX = CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_AMUX = CLBLM_L_X10Y136_SLICE_X13Y136_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_CMUX = CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_BMUX = CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_AMUX = CLBLM_L_X12Y124_SLICE_X16Y124_A5Q;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_BMUX = CLBLM_L_X12Y124_SLICE_X16Y124_B5Q;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A = CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B = CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C = CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_AMUX = CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_DMUX = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A = CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B = CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D = CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_AMUX = CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A = CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B = CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_AMUX = CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_BMUX = CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_CMUX = CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A = CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C = CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D = CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_BMUX = CLBLM_L_X12Y128_SLICE_X16Y128_BO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A = CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B = CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D = CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D = CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_AMUX = CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A = CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_BMUX = CLBLM_L_X12Y130_SLICE_X16Y130_B5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_AMUX = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_AMUX = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A = CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_CMUX = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_DMUX = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A = CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_AMUX = CLBLM_L_X12Y132_SLICE_X17Y132_AO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A = CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B = CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C = CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_CMUX = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_DMUX = CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C = CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_AMUX = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_BMUX = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_AMUX = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_BMUX = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_BMUX = CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B = CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_BMUX = CLBLM_R_X3Y127_SLICE_X2Y127_B5Q;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_CMUX = CLBLM_R_X3Y127_SLICE_X2Y127_C5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_AMUX = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B = CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C = CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D = CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C = CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D = CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_CMUX = CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B = CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A = CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C = CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_AMUX = CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_BMUX = CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D = CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_AMUX = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_CMUX = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A = CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_AMUX = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A = CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_BMUX = CLBLM_R_X3Y132_SLICE_X3Y132_B5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A = CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_BMUX = CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A = CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_BMUX = CLBLM_R_X5Y124_SLICE_X7Y124_B5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A = CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_DMUX = CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_BMUX = CLBLM_R_X5Y125_SLICE_X7Y125_B5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_CMUX = CLBLM_R_X5Y125_SLICE_X7Y125_C5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CMUX = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_AMUX = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_CMUX = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CMUX = CLBLM_R_X5Y127_SLICE_X6Y127_C5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_DMUX = CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_CMUX = CLBLM_R_X5Y127_SLICE_X7Y127_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A = CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B = CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CMUX = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_DMUX = CLBLM_R_X5Y128_SLICE_X6Y128_D5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A = CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B = CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_AMUX = CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_BMUX = CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CMUX = CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_DMUX = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_DMUX = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_AMUX = CLBLM_R_X5Y129_SLICE_X7Y129_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CMUX = CLBLM_R_X5Y129_SLICE_X7Y129_C5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_AMUX = CLBLM_R_X5Y130_SLICE_X6Y130_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_BMUX = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CMUX = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CMUX = CLBLM_R_X5Y130_SLICE_X7Y130_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A = CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_AMUX = CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CMUX = CLBLM_R_X5Y131_SLICE_X6Y131_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_DMUX = CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A = CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B = CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C = CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_AMUX = CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_BMUX = CLBLM_R_X5Y131_SLICE_X7Y131_B5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CMUX = CLBLM_R_X5Y131_SLICE_X7Y131_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_DMUX = CLBLM_R_X5Y131_SLICE_X7Y131_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_AMUX = CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_BMUX = CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CMUX = CLBLM_R_X5Y132_SLICE_X6Y132_C5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_DMUX = CLBLM_R_X5Y132_SLICE_X6Y132_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_AMUX = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_DMUX = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CMUX = CLBLM_R_X5Y133_SLICE_X6Y133_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_CMUX = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_DMUX = CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_AMUX = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A = CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B = CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_AMUX = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_BMUX = CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A = CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_AMUX = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_BMUX = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_CMUX = CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A = CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B = CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B = CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C = CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_AMUX = CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A = CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B = CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CMUX = CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A = CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B = CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CMUX = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A = CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B = CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_BMUX = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_BMUX = CLBLM_R_X7Y125_SLICE_X9Y125_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_DMUX = CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CMUX = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_AMUX = CLBLM_R_X7Y126_SLICE_X9Y126_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CMUX = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_DMUX = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_AMUX = CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_BMUX = CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_CMUX = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A = CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B = CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C = CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_AMUX = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_CMUX = CLBLM_R_X7Y128_SLICE_X8Y128_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_DMUX = CLBLM_R_X7Y128_SLICE_X8Y128_D5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A = CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_BMUX = CLBLM_R_X7Y128_SLICE_X9Y128_B5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_CMUX = CLBLM_R_X7Y128_SLICE_X9Y128_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_DMUX = CLBLM_R_X7Y128_SLICE_X9Y128_D5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_DMUX = CLBLM_R_X7Y129_SLICE_X8Y129_D5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_BMUX = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_CMUX = CLBLM_R_X7Y129_SLICE_X9Y129_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_BMUX = CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A = CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_BMUX = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CMUX = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_DMUX = CLBLM_R_X7Y130_SLICE_X9Y130_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CMUX = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_DMUX = CLBLM_R_X7Y131_SLICE_X8Y131_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_AMUX = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_BMUX = CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CMUX = CLBLM_R_X7Y131_SLICE_X9Y131_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_AMUX = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CMUX = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_AMUX = CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_BMUX = CLBLM_R_X7Y132_SLICE_X9Y132_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_CMUX = CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_BMUX = CLBLM_R_X7Y133_SLICE_X8Y133_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_DMUX = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A = CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_BMUX = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CMUX = CLBLM_R_X7Y133_SLICE_X9Y133_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_DMUX = CLBLM_R_X7Y133_SLICE_X9Y133_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B = CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C = CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_BMUX = CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A = CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B = CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_AMUX = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_BMUX = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_DMUX = CLBLM_R_X7Y134_SLICE_X9Y134_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_DMUX = CLBLM_R_X7Y135_SLICE_X8Y135_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A = CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B = CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_AMUX = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_BMUX = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_DMUX = CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A = CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_CMUX = CLBLM_R_X7Y136_SLICE_X8Y136_CO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_DMUX = CLBLM_R_X7Y136_SLICE_X9Y136_DO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B = CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A = CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_AMUX = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_BMUX = CLBLM_R_X11Y124_SLICE_X14Y124_B5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_BMUX = CLBLM_R_X11Y124_SLICE_X15Y124_B5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_CMUX = CLBLM_R_X11Y124_SLICE_X15Y124_C5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A = CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_AMUX = CLBLM_R_X11Y125_SLICE_X14Y125_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_BMUX = CLBLM_R_X11Y125_SLICE_X14Y125_B5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CMUX = CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_DMUX = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A = CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_AMUX = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A = CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_BMUX = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A = CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_AMUX = CLBLM_R_X11Y127_SLICE_X14Y127_A5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_BMUX = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_CMUX = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A = CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_BMUX = CLBLM_R_X11Y128_SLICE_X14Y128_B5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CMUX = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_DMUX = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A = CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_AMUX = CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A = CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B = CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_DMUX = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_AMUX = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_DMUX = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A = CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_AMUX = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_AMUX = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_BMUX = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CMUX = CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_DMUX = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A = CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_BMUX = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_AMUX = CLBLM_R_X11Y132_SLICE_X15Y132_A5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_BMUX = CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_CMUX = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CMUX = CLBLM_R_X11Y133_SLICE_X14Y133_C5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_DMUX = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_DMUX = CLBLM_R_X11Y133_SLICE_X15Y133_D5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_BMUX = CLBLM_R_X11Y134_SLICE_X14Y134_B5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CMUX = CLBLM_R_X11Y134_SLICE_X14Y134_C5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_DMUX = CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_AMUX = CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_CMUX = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_AMUX = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_AMUX = CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B = CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C = CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A = CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B = CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C = CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D = CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_AMUX = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_BMUX = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D = CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B = CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_AMUX = CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B = CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_CMUX = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_AMUX = CLBLM_R_X13Y129_SLICE_X18Y129_AO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_CMUX = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A = CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A = CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_BMUX = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_DMUX = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D = CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_AMUX = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_CMUX = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A = CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B = CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D = CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_AMUX = CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_BMUX = CLBLM_R_X13Y131_SLICE_X18Y131_BO5;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B = CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C = CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D = CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D = CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_AMUX = CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_BMUX = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A = CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B = CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C = CLBLM_R_X13Y133_SLICE_X18Y133_CO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D = CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_AMUX = CLBLM_R_X13Y133_SLICE_X18Y133_AO5;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_BMUX = CLBLM_R_X13Y133_SLICE_X18Y133_BO5;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A = CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B = CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D = CLBLM_R_X13Y133_SLICE_X19Y133_DO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_AMUX = CLBLM_R_X13Y133_SLICE_X19Y133_AO5;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_BMUX = CLBLM_R_X13Y133_SLICE_X19Y133_BO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_AMUX = CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A = CLBLM_R_X13Y134_SLICE_X19Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B = CLBLM_R_X13Y134_SLICE_X19Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C = CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D = CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A = CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B = CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C = CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D = CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B = CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C = CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D = CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_OQ = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_TQ = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X4Y125_SLICE_X5Y125_CQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X4Y126_SLICE_X5Y126_CQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X11Y124_SLICE_X15Y124_B5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X7Y131_SLICE_X9Y131_C5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_L_X10Y125_SLICE_X13Y125_A5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ = CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X5Y133_SLICE_X6Y133_C5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X8Y132_SLICE_X11Y132_C5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y133_SLICE_X19Y133_BO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X13Y133_SLICE_X19Y133_AO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A2 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A4 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B5 = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B6 = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C1 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C2 = CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C5 = CLBLM_R_X5Y131_SLICE_X6Y131_C5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D2 = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D3 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D5 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D6 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A3 = CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A4 = CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A5 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B1 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B3 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B4 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B5 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B6 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C3 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C4 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C5 = CLBLM_R_X5Y132_SLICE_X6Y132_C5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C6 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D2 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D3 = CLBLM_R_X7Y129_SLICE_X8Y129_D5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D5 = CLBLM_R_X11Y124_SLICE_X15Y124_B5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_O = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y152_O = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign LIOB33_X0Y151_IOB_X0Y151_O = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = CLBLM_R_X3Y127_SLICE_X2Y127_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = CLBLM_L_X8Y134_SLICE_X10Y134_D5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = CLBLM_R_X5Y130_SLICE_X7Y130_C5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = CLBLM_R_X7Y130_SLICE_X9Y130_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = CLBLM_L_X8Y129_SLICE_X11Y129_DQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign LIOB33_X0Y153_IOB_X0Y154_O = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign LIOB33_X0Y153_IOB_X0Y153_O = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A2 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A3 = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B3 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B4 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B5 = CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C1 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C2 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C3 = CLBLL_L_X4Y125_SLICE_X5Y125_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C5 = CLBLM_R_X5Y131_SLICE_X7Y131_B5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D2 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D5 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A1 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A2 = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A5 = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B1 = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B2 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B4 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C1 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C2 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C4 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C5 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D1 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D3 = CLBLM_R_X5Y132_SLICE_X7Y132_DQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D5 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign LIOB33_X0Y155_IOB_X0Y155_O = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X13Y133_SLICE_X19Y133_AO5;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A1 = CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A4 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A5 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B2 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B4 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B5 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B6 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C1 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C2 = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C5 = CLBLM_R_X5Y131_SLICE_X7Y131_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C6 = CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D3 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D4 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D5 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A2 = CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A3 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_DQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A5 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A6 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_AX = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B2 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B3 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B4 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B5 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B6 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_BX = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C3 = CLBLM_R_X5Y132_SLICE_X6Y132_DQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C4 = CLBLM_L_X8Y129_SLICE_X10Y129_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C5 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D1 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D2 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D5 = CLBLM_R_X5Y127_SLICE_X7Y127_DQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D6 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D4 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A1 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A2 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A3 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A5 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A6 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B1 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B2 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B4 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B6 = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C5 = CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C1 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C3 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A1 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A3 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A4 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A5 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A6 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B1 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B2 = CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B3 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B4 = CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B5 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C1 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C2 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C6 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D2 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D1 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = CLBLL_L_X2Y123_SLICE_X1Y123_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = CLBLM_R_X3Y124_SLICE_X2Y124_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D3 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D4 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D5 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X4Y125_SLICE_X5Y125_CQ;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A1 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A2 = CLBLM_R_X5Y133_SLICE_X6Y133_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A3 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A5 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B1 = CLBLM_R_X5Y131_SLICE_X7Y131_B5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B3 = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B5 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B6 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C1 = CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D1 = CLBLM_R_X5Y127_SLICE_X7Y127_C5Q;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A1 = CLBLL_L_X4Y129_SLICE_X4Y129_DQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A3 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A4 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A5 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A6 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B2 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B3 = CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A2 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A3 = CLBLM_R_X3Y124_SLICE_X2Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A4 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A5 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B1 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B2 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B3 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B4 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C2 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C3 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C6 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D6 = 1'b1;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A6 = CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B3 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B4 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B5 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B6 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C2 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C4 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C5 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C6 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A1 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A3 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A4 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A6 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign LIOB33_X0Y163_IOB_X0Y163_O = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_AX = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B1 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B5 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A1 = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A4 = CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A5 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A6 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C1 = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B3 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B4 = CLBLM_R_X3Y127_SLICE_X2Y127_BQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B6 = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D1 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D2 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A1 = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A2 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A3 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_DQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B1 = CLBLL_L_X4Y132_SLICE_X4Y132_DQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B2 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B3 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C1 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C2 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D1 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D3 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D4 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D6 = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A2 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A3 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A4 = CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B4 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X4Y126_SLICE_X5Y126_CQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A1 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A2 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A4 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A5 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B1 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B2 = CLBLL_L_X4Y126_SLICE_X5Y126_A5Q;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B3 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B4 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B5 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C1 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_C5Q;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C3 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C4 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C5 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C6 = CLBLM_R_X7Y129_SLICE_X8Y129_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B2 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B3 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_AX = CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D2 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D3 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D4 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D1 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D2 = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D3 = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A1 = CLBLM_R_X7Y126_SLICE_X9Y126_DQ;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A2 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A5 = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B2 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B4 = CLBLM_L_X8Y127_SLICE_X10Y127_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C5 = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A1 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A3 = CLBLM_L_X8Y127_SLICE_X11Y127_D5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A4 = CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B1 = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B3 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B4 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_D5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B6 = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C1 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C2 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C3 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C5 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C6 = CLBLM_R_X5Y127_SLICE_X6Y127_C5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D1 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D2 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D3 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D5 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D6 = CLBLM_R_X5Y127_SLICE_X6Y127_C5Q;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A1 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A3 = CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A4 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A5 = CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A6 = CLBLL_L_X2Y123_SLICE_X1Y123_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B2 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B3 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B5 = CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C2 = CLBLM_R_X3Y127_SLICE_X2Y127_CQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C3 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C4 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C5 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C6 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D2 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D3 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A4 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A5 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B1 = CLBLL_L_X4Y129_SLICE_X4Y129_DQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B2 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B5 = CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A1 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A2 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_C5Q;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A4 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A5 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A6 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_AX = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B1 = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B2 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B4 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B5 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B6 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C3 = CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C4 = CLBLM_L_X10Y136_SLICE_X13Y136_A5Q;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C5 = CLBLL_L_X4Y129_SLICE_X5Y129_C5Q;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D3 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D5 = CLBLM_L_X8Y129_SLICE_X11Y129_C5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X8Y132_SLICE_X11Y132_C5Q;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D3 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign LIOB33_X0Y171_IOB_X0Y172_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y171_IOB_X0Y171_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D5 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A6 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A2 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A3 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A4 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_D5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B1 = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B2 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B3 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B4 = CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B5 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C2 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C3 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C4 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C5 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C6 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C5 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C6 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D2 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D3 = CLBLM_R_X3Y129_SLICE_X3Y129_DQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D5 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A1 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A4 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A5 = CLBLM_R_X3Y127_SLICE_X2Y127_C5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A6 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A3 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B1 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B2 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B4 = CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B6 = CLBLM_L_X10Y125_SLICE_X12Y125_B5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C1 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C2 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C3 = CLBLM_R_X3Y129_SLICE_X2Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C4 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D1 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D1 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D2 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D4 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D5 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A4 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D4 = CLBLM_R_X7Y133_SLICE_X8Y133_B5Q;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D5 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D6 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C4 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D4 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A1 = CLBLM_L_X12Y124_SLICE_X16Y124_B5Q;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A2 = CLBLM_L_X12Y124_SLICE_X16Y124_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A3 = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A4 = CLBLM_L_X12Y124_SLICE_X16Y124_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A5 = CLBLM_L_X12Y124_SLICE_X16Y124_A5Q;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B3 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y173_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y173_IOB_X0Y174_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A1 = CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B1 = CLBLM_L_X12Y124_SLICE_X16Y124_B5Q;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B2 = CLBLM_L_X12Y124_SLICE_X16Y124_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B3 = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B4 = CLBLM_L_X12Y124_SLICE_X16Y124_CQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B5 = CLBLM_L_X12Y124_SLICE_X16Y124_A5Q;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A3 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C2 = CLBLM_L_X12Y124_SLICE_X16Y124_CQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A4 = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C4 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C5 = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A6 = CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D4 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B3 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B4 = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B5 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B6 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C1 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C3 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C4 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C5 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C6 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A1 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A3 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A4 = CLBLM_L_X8Y129_SLICE_X10Y129_D5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A6 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D1 = CLBLM_L_X8Y132_SLICE_X11Y132_C5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D2 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D3 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D4 = CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D5 = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A1 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A3 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A5 = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_AX = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B3 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B4 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B5 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A2 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A3 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A4 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A5 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B2 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B3 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B4 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B5 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B6 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C2 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C3 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C4 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C5 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C6 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D2 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D3 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D4 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D5 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A1 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A4 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A5 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B2 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B3 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B4 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B6 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C1 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C3 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C4 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C6 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D1 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D4 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D5 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D6 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B5 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X5Y133_SLICE_X6Y133_C5Q;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A1 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A2 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A3 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A5 = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B1 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B2 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B3 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B4 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B6 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C1 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C2 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C3 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C4 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C5 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C6 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A1 = CLBLL_L_X4Y125_SLICE_X5Y125_C5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A3 = CLBLM_R_X3Y127_SLICE_X2Y127_C5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B6 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C6 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C1 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C2 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A3 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A4 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C3 = CLBLM_L_X8Y126_SLICE_X11Y126_DQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B1 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C4 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B3 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B4 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B6 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C1 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C4 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C6 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D1 = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D2 = CLBLM_R_X5Y128_SLICE_X7Y128_DQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D3 = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D4 = CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D5 = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D6 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D3 = CLBLM_R_X7Y135_SLICE_X8Y135_D5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D4 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A1 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A4 = CLBLM_L_X12Y130_SLICE_X16Y130_B5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A6 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B1 = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B2 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B5 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B6 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C1 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C2 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C3 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C4 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C6 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D2 = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D3 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D4 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D5 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D6 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D5 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B4 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B5 = CLBLM_R_X7Y132_SLICE_X9Y132_B5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B6 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A1 = CLBLM_R_X3Y129_SLICE_X3Y129_DQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A2 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A3 = CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A4 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A5 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B2 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B4 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B5 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C1 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C2 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C3 = CLBLM_R_X7Y132_SLICE_X9Y132_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C4 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C6 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D1 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D2 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D3 = CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D5 = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D6 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A1 = CLBLM_R_X3Y129_SLICE_X3Y129_DQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A4 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A5 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A6 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A1 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A2 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A3 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B1 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B2 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B3 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C2 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C3 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C4 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D1 = CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D2 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D3 = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D4 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D5 = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D6 = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A1 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A2 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A3 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A4 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A5 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B1 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B2 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B3 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B5 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C1 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C2 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C6 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D2 = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D3 = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D4 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D5 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A1 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A3 = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A4 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A5 = CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A6 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B2 = CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B3 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B4 = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B5 = CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B6 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C1 = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C2 = CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C3 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C4 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C5 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C6 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D1 = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D2 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D3 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D6 = CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A1 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A2 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A3 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A4 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A6 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B1 = CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B3 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B4 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B5 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C1 = CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C1 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C3 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C4 = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C5 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C6 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C2 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D2 = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D3 = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D4 = CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D5 = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D6 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign LIOB33_X0Y63_IOB_X0Y64_O = CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D3 = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign RIOB33_X105Y151_IOB_X1Y152_O = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y151_O = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C1 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C2 = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A1 = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A2 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A3 = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A4 = CLBLL_L_X4Y128_SLICE_X5Y128_CQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A5 = CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C1 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C2 = CLBLM_R_X11Y133_SLICE_X15Y133_D5Q;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B1 = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B2 = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B3 = CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B4 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B5 = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B6 = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C1 = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C2 = CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C3 = CLBLL_L_X4Y128_SLICE_X4Y128_C5Q;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C4 = CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C5 = CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C6 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D1 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D2 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D3 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D4 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D5 = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D6 = CLBLM_R_X13Y129_SLICE_X18Y129_AO5;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A1 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A3 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A4 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A5 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A6 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B1 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B2 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B3 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B5 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B6 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A1 = CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C1 = CLBLM_L_X8Y125_SLICE_X10Y125_C5Q;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C2 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A2 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C6 = CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C3 = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A3 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A5 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D2 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D3 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D4 = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A6 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D5 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D6 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign LIOB33_X0Y65_IOB_X0Y65_O = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign LIOB33_X0Y65_IOB_X0Y66_O = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign RIOB33_X105Y153_IOB_X1Y154_O = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_O = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign LIOB33_X0Y159_IOB_X0Y159_O = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D5 = CLBLM_R_X7Y135_SLICE_X9Y135_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A1 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A2 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A3 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B1 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B2 = CLBLM_L_X8Y130_SLICE_X11Y130_D5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B3 = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B4 = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B5 = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B6 = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C1 = CLBLM_R_X3Y130_SLICE_X3Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C2 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C3 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C4 = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C5 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C6 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D2 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D3 = CLBLM_L_X8Y130_SLICE_X11Y130_D5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D4 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D5 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D6 = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X11Y124_SLICE_X15Y124_B5Q;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A1 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A5 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A6 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B5 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C1 = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C2 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C3 = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C4 = CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C5 = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C6 = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_C5Q;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D1 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D4 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D5 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y155_O = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_O = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign LIOB33_X0Y187_IOB_X0Y187_O = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A4 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B1 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B2 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C2 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C3 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C4 = CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A1 = CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A2 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A3 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A4 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A5 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A6 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_AX = CLBLM_R_X13Y131_SLICE_X18Y131_BO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B1 = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C2 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B2 = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B3 = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B4 = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B5 = CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C3 = CLBLM_L_X8Y127_SLICE_X11Y127_DQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B6 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C4 = CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C2 = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C3 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C5 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C6 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D1 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D2 = CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D3 = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D4 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D5 = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D6 = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A1 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A2 = CLBLM_L_X8Y128_SLICE_X10Y128_D5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A3 = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A4 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A5 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A6 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_AX = CLBLL_L_X4Y129_SLICE_X4Y129_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B1 = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B2 = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B3 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B4 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B6 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D6 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y157_O = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C2 = CLBLM_L_X12Y132_SLICE_X17Y132_AO5;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C3 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C4 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C5 = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C6 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D1 = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D2 = CLBLM_L_X8Y130_SLICE_X11Y130_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D2 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D3 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D4 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D5 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D4 = CLBLM_R_X5Y124_SLICE_X7Y124_B5Q;
  assign LIOB33_X0Y189_IOB_X0Y190_O = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign LIOB33_X0Y189_IOB_X0Y189_O = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign LIOB33_X0Y161_IOB_X0Y162_O = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y161_IOB_X0Y161_O = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B2 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B3 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C4 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A2 = CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A3 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A4 = CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A5 = CLBLM_R_X11Y133_SLICE_X14Y133_C5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_AX = CLBLM_R_X11Y132_SLICE_X15Y132_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B1 = CLBLM_L_X10Y132_SLICE_X12Y132_DQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B2 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B3 = CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B4 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B6 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C2 = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C3 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C4 = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C5 = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D1 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D3 = CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D4 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D6 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign RIOB33_X105Y159_IOB_X1Y159_O = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A1 = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A2 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A3 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A4 = CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B1 = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B4 = CLBLM_L_X8Y128_SLICE_X10Y128_D5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B5 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C1 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C2 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C3 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C4 = CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C5 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D1 = CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D2 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D4 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D5 = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y191_O = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign LIOB33_X0Y191_IOB_X0Y192_O = CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X8Y132_SLICE_X11Y132_C5Q;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_L_X10Y125_SLICE_X13Y125_A5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A3 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A4 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A5 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A6 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C4 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D1 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D2 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D3 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D4 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D5 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A1 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A2 = CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A3 = CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A4 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A5 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D6 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_AX = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B1 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B2 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B3 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B5 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B6 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_BX = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C4 = CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C6 = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D1 = CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D6 = CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A1 = CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A3 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A5 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A6 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B2 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B3 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B4 = CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C4 = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C5 = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D1 = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A2 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A3 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A4 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A6 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B2 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B3 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B5 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B6 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C1 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C2 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C5 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C6 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A4 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A5 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B2 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B5 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B6 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C1 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C2 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C3 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C4 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C6 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A2 = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D1 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D2 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D3 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D4 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A5 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D6 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A6 = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C3 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C5 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B2 = 1'b1;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A3 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A4 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A5 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D1 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B2 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B3 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B5 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B6 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C1 = CLBLM_L_X10Y132_SLICE_X13Y132_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C2 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C4 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C5 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C6 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A1 = CLBLM_L_X8Y127_SLICE_X10Y127_D5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A3 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A4 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A5 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D4 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D1 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D3 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D5 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D6 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B3 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B4 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D6 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A1 = CLBLM_L_X8Y128_SLICE_X11Y128_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A3 = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A4 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A1 = CLBLM_L_X8Y132_SLICE_X11Y132_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A4 = CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A6 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B1 = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B2 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_DQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B6 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C1 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C2 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C3 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A5 = CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A6 = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D2 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_AX = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B1 = CLBLM_L_X8Y134_SLICE_X10Y134_C5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B2 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B3 = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B4 = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A3 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A5 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A6 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B1 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B6 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B3 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B4 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B6 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C1 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C2 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C3 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C6 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D1 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D2 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D3 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C2 = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A1 = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A2 = CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A3 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A4 = CLBLM_L_X10Y126_SLICE_X12Y126_C5Q;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A5 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C4 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_AX = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B1 = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B2 = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C5 = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B4 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B5 = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B6 = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C1 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C2 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C3 = CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C4 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C5 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C6 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D1 = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D2 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D3 = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D4 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D5 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D6 = CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign RIOB33_X105Y165_IOB_X1Y165_O = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D1 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D2 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D5 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y197_O = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A1 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A3 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A4 = CLBLM_L_X10Y127_SLICE_X12Y127_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B1 = CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B2 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B3 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B5 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C2 = CLBLM_L_X10Y127_SLICE_X12Y127_D5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C3 = CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C4 = CLBLM_L_X10Y125_SLICE_X12Y125_CQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C5 = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D1 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D3 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D4 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D5 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A1 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A3 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A5 = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B2 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B3 = CLBLM_L_X10Y125_SLICE_X12Y125_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B4 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C4 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C5 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C6 = CLBLM_L_X10Y127_SLICE_X12Y127_D5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D2 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D3 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D4 = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D6 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C4 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C5 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C6 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A1 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A2 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A3 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A5 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B1 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B2 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B3 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B5 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C1 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C2 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C3 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C5 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D1 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D2 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D3 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D5 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A2 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D2 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A3 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A4 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B1 = CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B2 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B3 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B4 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B5 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D5 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C1 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C2 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C3 = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C4 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C5 = CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C6 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign RIOB33_X105Y167_IOB_X1Y167_O = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D1 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D2 = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D3 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D4 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D5 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D6 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C4 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B5 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A1 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A2 = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A3 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A4 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A5 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A6 = CLBLM_R_X7Y128_SLICE_X9Y128_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_AX = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B2 = CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B3 = CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B4 = CLBLM_L_X8Y134_SLICE_X11Y134_D5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B5 = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B6 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C1 = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C2 = CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C3 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C4 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C5 = CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C6 = CLBLM_R_X7Y130_SLICE_X9Y130_D5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D1 = CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D2 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D6 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C4 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A1 = CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A3 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A6 = CLBLM_L_X10Y128_SLICE_X13Y128_A5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D5 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C6 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B1 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B2 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B3 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B4 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C2 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C3 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C5 = CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X5Y133_SLICE_X6Y133_C5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D1 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D3 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D4 = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D5 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A5 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A3 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A4 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A5 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A6 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B1 = CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B2 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B3 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B5 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B6 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C1 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C2 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C3 = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C4 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C5 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C6 = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D2 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D4 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B4 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B5 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A1 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A2 = CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A3 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A4 = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A5 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A6 = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B1 = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B2 = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B3 = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B4 = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B5 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B6 = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C2 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C3 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C4 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C6 = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D2 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D3 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D4 = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D6 = CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C4 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A2 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A3 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A4 = CLBLL_L_X4Y128_SLICE_X5Y128_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A5 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A6 = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B1 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B2 = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B3 = CLBLM_R_X5Y125_SLICE_X7Y125_C5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B4 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B5 = CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B6 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C1 = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C2 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C3 = CLBLM_L_X10Y129_SLICE_X12Y129_B5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C4 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C5 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C6 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D2 = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D5 = CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D6 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A3 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A4 = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_C5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B1 = CLBLM_R_X11Y127_SLICE_X14Y127_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B2 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B5 = CLBLM_L_X8Y127_SLICE_X11Y127_C5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C2 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C4 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C6 = CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D2 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D3 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D4 = CLBLM_L_X8Y134_SLICE_X10Y134_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D5 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A2 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A3 = CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B6 = CLBLM_L_X10Y125_SLICE_X13Y125_A5Q;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A4 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A6 = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B2 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B3 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B4 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C2 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C3 = CLBLM_R_X13Y133_SLICE_X18Y133_BO5;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C4 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C5 = CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C6 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D2 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D3 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D4 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D5 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A2 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A3 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A4 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A5 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B1 = CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B2 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B4 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B5 = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C1 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C2 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C3 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C4 = CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C6 = CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D1 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D2 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D3 = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D4 = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D5 = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D6 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A3 = CLBLM_R_X11Y125_SLICE_X14Y125_B5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A1 = CLBLM_R_X7Y128_SLICE_X9Y128_D5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A2 = CLBLM_R_X7Y129_SLICE_X8Y129_D5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B1 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B4 = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B5 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B6 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_BX = CLBLM_L_X12Y128_SLICE_X16Y128_BO5;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C1 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C2 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C4 = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C6 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D3 = CLBLM_R_X11Y128_SLICE_X14Y128_B5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D5 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D6 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C4 = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A2 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A4 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A5 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A6 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_AX = CLBLM_L_X8Y129_SLICE_X10Y129_DQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B1 = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B2 = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B3 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B4 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B5 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B6 = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C5 = CLBLM_L_X10Y125_SLICE_X13Y125_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A1 = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C1 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C2 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C4 = CLBLM_L_X10Y126_SLICE_X12Y126_C5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C5 = CLBLM_L_X10Y129_SLICE_X13Y129_CQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C6 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B5 = CLBLL_L_X4Y126_SLICE_X5Y126_C5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B6 = CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B1 = CLBLM_R_X3Y127_SLICE_X2Y127_B5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D3 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D4 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D5 = CLBLM_R_X11Y132_SLICE_X15Y132_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D6 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D5 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A1 = CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A2 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A4 = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B1 = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B2 = CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B3 = CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C1 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C3 = CLBLM_R_X13Y133_SLICE_X18Y133_BO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C4 = CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C5 = CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D1 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D5 = CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A1 = CLBLM_R_X13Y133_SLICE_X18Y133_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A2 = CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A3 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A4 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A5 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A6 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B1 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B2 = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B4 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B5 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C1 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C2 = CLBLM_R_X13Y133_SLICE_X18Y133_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C3 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C4 = CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C5 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D1 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D3 = CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D4 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D6 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A2 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A5 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A1 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A3 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B5 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A5 = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A6 = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C3 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C5 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B5 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C1 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D5 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C5 = CLBLM_R_X7Y135_SLICE_X9Y135_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D1 = CLBLM_L_X10Y129_SLICE_X13Y129_C5Q;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D2 = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D5 = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D6 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A1 = CLBLM_L_X10Y129_SLICE_X12Y129_B5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A2 = CLBLM_L_X10Y128_SLICE_X13Y128_A5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A3 = CLBLM_L_X8Y132_SLICE_X11Y132_C5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B2 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B3 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A3 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A6 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_AX = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A1 = CLBLL_L_X4Y125_SLICE_X5Y125_BO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B1 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B2 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C4 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B5 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C1 = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C2 = CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C4 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C5 = CLBLL_L_X4Y125_SLICE_X5Y125_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D1 = CLBLM_R_X11Y133_SLICE_X14Y133_DQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D5 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D2 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D3 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D4 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D5 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A1 = CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A3 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A4 = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B2 = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B3 = CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B5 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A3 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A4 = CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A5 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B1 = CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B3 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B4 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B5 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_T1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C1 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C3 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D3 = CLBLM_R_X11Y132_SLICE_X15Y132_B5Q;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D6 = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A5 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C5 = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C6 = CLBLM_R_X11Y133_SLICE_X15Y133_D5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A2 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A4 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A5 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_AX = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B1 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B2 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B4 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B5 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C2 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C3 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C4 = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C5 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C6 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = CLBLM_L_X8Y133_SLICE_X10Y133_D5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = CLBLM_R_X7Y133_SLICE_X8Y133_DQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A1 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A2 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A3 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A5 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A6 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_AX = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B1 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B2 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B3 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B6 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = CLBLM_R_X7Y129_SLICE_X9Y129_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C1 = CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C2 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C5 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D1 = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D2 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D3 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D4 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D5 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D6 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = CLBLM_R_X5Y129_SLICE_X7Y129_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C1 = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C5 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A1 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A4 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C6 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B1 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A1 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A2 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A4 = CLBLM_R_X11Y124_SLICE_X14Y124_B5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A5 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A6 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B6 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B4 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B5 = CLBLM_R_X11Y124_SLICE_X15Y124_C5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D1 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C2 = CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C5 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A2 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A3 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A4 = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D3 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D5 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B1 = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B2 = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B3 = CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A2 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C5 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B3 = CLBLM_R_X11Y124_SLICE_X15Y124_C5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B4 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B5 = CLBLL_L_X4Y130_SLICE_X4Y130_C5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D3 = CLBLM_R_X11Y133_SLICE_X14Y133_C5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D4 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D6 = CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A1 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A2 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A4 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A5 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B2 = CLBLL_L_X4Y127_SLICE_X4Y127_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B3 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_C5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C5 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = CLBLM_R_X11Y131_SLICE_X14Y131_DQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_C5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D2 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D4 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = CLBLM_L_X8Y129_SLICE_X10Y129_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = CLBLL_L_X4Y132_SLICE_X4Y132_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = CLBLM_L_X8Y130_SLICE_X10Y130_D5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A2 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A3 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A4 = CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A5 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A6 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = CLBLM_L_X12Y130_SLICE_X16Y130_B5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B2 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B4 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B5 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B6 = CLBLM_R_X5Y129_SLICE_X7Y129_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C2 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C3 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C5 = CLBLL_L_X4Y127_SLICE_X4Y127_DQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D1 = CLBLL_L_X4Y126_SLICE_X5Y126_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D2 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D3 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D5 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D6 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A2 = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A3 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A4 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A5 = CLBLM_R_X11Y132_SLICE_X15Y132_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A6 = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B1 = CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B2 = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B5 = CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B6 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C2 = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C3 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C4 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C5 = CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C6 = CLBLM_R_X5Y132_SLICE_X7Y132_DQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D1 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D2 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D3 = CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D4 = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D6 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A2 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A3 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A5 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B1 = CLBLL_L_X4Y127_SLICE_X4Y127_D5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B3 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B4 = CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B5 = CLBLM_R_X11Y125_SLICE_X14Y125_C5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C1 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C3 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C5 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D1 = CLBLM_R_X5Y132_SLICE_X6Y132_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D2 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D3 = CLBLL_L_X4Y128_SLICE_X5Y128_C5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D5 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D6 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A3 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A4 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A5 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A6 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B1 = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B2 = CLBLM_R_X3Y126_SLICE_X3Y126_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B3 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B4 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B6 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C3 = CLBLM_R_X3Y132_SLICE_X3Y132_B5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C4 = CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C5 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = CLBLM_L_X10Y136_SLICE_X13Y136_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = CLBLM_L_X8Y133_SLICE_X10Y133_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_AX = CLBLM_L_X10Y133_SLICE_X13Y133_CQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = CLBLM_L_X8Y129_SLICE_X10Y129_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = CLBLM_R_X5Y132_SLICE_X7Y132_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_BX = CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = CLBLM_L_X10Y133_SLICE_X12Y133_DQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A2 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A3 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A6 = CLBLM_R_X7Y128_SLICE_X9Y128_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = CLBLM_L_X8Y129_SLICE_X11Y129_D5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B1 = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B5 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C4 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C6 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D2 = CLBLL_L_X4Y127_SLICE_X4Y127_DQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = CLBLM_L_X10Y132_SLICE_X12Y132_DQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D3 = CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D5 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A1 = CLBLM_R_X11Y124_SLICE_X14Y124_B5Q;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A2 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A3 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A4 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B2 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B3 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B4 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C1 = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C2 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C3 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C4 = CLBLM_R_X5Y129_SLICE_X7Y129_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C5 = CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C6 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D1 = CLBLM_L_X10Y125_SLICE_X12Y125_B5Q;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D2 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D3 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D4 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D5 = CLBLM_L_X10Y126_SLICE_X12Y126_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A2 = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A3 = CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A4 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_AX = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B2 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B3 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B4 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B6 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C1 = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C2 = CLBLM_R_X5Y125_SLICE_X7Y125_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C3 = CLBLM_L_X8Y128_SLICE_X10Y128_DQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C4 = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C5 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C6 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D1 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D2 = CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D3 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D5 = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D6 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign RIOB33_X105Y183_IOB_X1Y183_O = 1'b0;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A2 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A3 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A6 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B1 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B4 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B5 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B6 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C1 = CLBLL_L_X4Y127_SLICE_X4Y127_C5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C2 = CLBLL_L_X4Y129_SLICE_X4Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C4 = CLBLL_L_X4Y129_SLICE_X5Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C5 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C6 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A1 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A4 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A5 = CLBLM_L_X10Y133_SLICE_X13Y133_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D1 = CLBLL_L_X4Y129_SLICE_X4Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D2 = CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D3 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D4 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D6 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A6 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B1 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B2 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B3 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B5 = CLBLM_R_X11Y134_SLICE_X14Y134_C5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C1 = CLBLM_L_X8Y129_SLICE_X11Y129_D5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C2 = CLBLM_L_X10Y133_SLICE_X13Y133_CQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C3 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C4 = CLBLM_R_X7Y134_SLICE_X9Y134_D5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C6 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D2 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D3 = CLBLM_L_X10Y133_SLICE_X13Y133_DQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A1 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A2 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A4 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A6 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D4 = CLBLM_R_X11Y132_SLICE_X15Y132_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D5 = CLBLM_R_X7Y133_SLICE_X9Y133_C5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A2 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A4 = CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A5 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B1 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B2 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B4 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B1 = CLBLM_L_X8Y133_SLICE_X10Y133_B5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B6 = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C1 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C2 = CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C3 = CLBLM_R_X11Y128_SLICE_X14Y128_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A1 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A4 = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A5 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D2 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D4 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D5 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B1 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B5 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D3 = CLBLM_L_X10Y133_SLICE_X12Y133_DQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D4 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A1 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A3 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A4 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A5 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A6 = CLBLM_R_X11Y124_SLICE_X15Y124_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B1 = CLBLM_R_X11Y128_SLICE_X14Y128_B5Q;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B2 = CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B3 = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B4 = CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B5 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B6 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C1 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C2 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C3 = CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C5 = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C6 = CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D1 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D3 = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D4 = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D5 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D6 = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A1 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A2 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A3 = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A5 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B3 = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B4 = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B5 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B6 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y133_SLICE_X19Y133_BO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C3 = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C4 = CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C5 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C6 = CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D1 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D2 = CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D3 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D5 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B3 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D6 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A2 = CLBLM_R_X3Y132_SLICE_X3Y132_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A3 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A4 = CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A6 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B2 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B3 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B4 = CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B6 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C2 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C4 = CLBLM_R_X5Y129_SLICE_X7Y129_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C5 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A1 = CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D1 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D2 = CLBLM_R_X5Y130_SLICE_X6Y130_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D4 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D5 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A3 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A5 = CLBLM_R_X11Y128_SLICE_X14Y128_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B1 = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B3 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B4 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B5 = CLBLM_R_X11Y134_SLICE_X14Y134_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B6 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A4 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A5 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C1 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C2 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C3 = CLBLM_R_X7Y133_SLICE_X8Y133_B5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B2 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B3 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B4 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B5 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A1 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A2 = CLBLM_R_X5Y131_SLICE_X6Y131_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A3 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A4 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C3 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C4 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C5 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C6 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B1 = CLBLM_R_X5Y131_SLICE_X7Y131_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B2 = CLBLM_R_X3Y130_SLICE_X2Y130_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D2 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B5 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B2 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C2 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C3 = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D5 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C5 = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A4 = CLBLM_R_X7Y128_SLICE_X8Y128_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A1 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A2 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D2 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D3 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D4 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D5 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B2 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B3 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B5 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B6 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C1 = CLBLM_L_X10Y129_SLICE_X13Y129_C5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C2 = CLBLM_L_X8Y124_SLICE_X10Y124_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C3 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C4 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C5 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D6 = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D2 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D3 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D4 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D5 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D6 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C2 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A1 = CLBLM_R_X3Y127_SLICE_X2Y127_B5Q;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A2 = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A4 = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A5 = CLBLM_L_X8Y129_SLICE_X10Y129_DQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B1 = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B2 = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B3 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B4 = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B5 = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B6 = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C1 = CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C2 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C4 = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C5 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C6 = CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X4Y125_SLICE_X5Y125_CQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D2 = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D4 = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D6 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A2 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A5 = CLBLM_L_X8Y129_SLICE_X11Y129_C5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A6 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B1 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B2 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B5 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B6 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C2 = CLBLM_L_X10Y126_SLICE_X12Y126_DQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A2 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C5 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D1 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D5 = CLBLM_R_X5Y128_SLICE_X7Y128_DQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D6 = CLBLM_R_X5Y129_SLICE_X7Y129_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A1 = CLBLM_R_X11Y131_SLICE_X14Y131_DQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A2 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A3 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A5 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B1 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B3 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B4 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C1 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C2 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C3 = CLBLL_L_X4Y131_SLICE_X4Y131_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C4 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C6 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D4 = CLBLL_L_X4Y130_SLICE_X4Y130_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D6 = CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A1 = CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A2 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A3 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A4 = CLBLM_L_X10Y127_SLICE_X12Y127_D5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A5 = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_AX = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B2 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B3 = CLBLM_R_X11Y133_SLICE_X14Y133_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B6 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A1 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A2 = CLBLM_R_X7Y128_SLICE_X9Y128_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C3 = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C4 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A5 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A6 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_AX = CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D1 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D2 = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D3 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D4 = CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D5 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A3 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B5 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C3 = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C4 = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C6 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B6 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C2 = CLBLL_L_X4Y131_SLICE_X5Y131_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B4 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B5 = CLBLM_R_X11Y134_SLICE_X14Y134_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B6 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D3 = CLBLM_R_X5Y133_SLICE_X6Y133_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C1 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C4 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C6 = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D4 = CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B1 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B3 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D1 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D2 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D3 = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D6 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C2 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C3 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C5 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D1 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D3 = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D4 = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D5 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D6 = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C3 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_DQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C5 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X4Y126_SLICE_X5Y126_CQ;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A1 = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A2 = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A3 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A4 = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A5 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A6 = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B1 = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B2 = CLBLM_R_X11Y125_SLICE_X14Y125_A5Q;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B3 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B4 = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B5 = CLBLM_R_X11Y127_SLICE_X14Y127_A5Q;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B6 = CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C1 = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C2 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C3 = CLBLM_L_X8Y128_SLICE_X11Y128_C5Q;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C4 = CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C5 = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C6 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D2 = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D3 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D5 = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D6 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y133_SLICE_X19Y133_BO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D1 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A2 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A3 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A5 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A6 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C3 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B1 = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B2 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B3 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B4 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B5 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B6 = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D5 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C4 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C5 = CLBLM_R_X7Y134_SLICE_X9Y134_D5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C1 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C2 = CLBLL_L_X4Y130_SLICE_X4Y130_C5Q;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C3 = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C4 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C5 = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C6 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D2 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D3 = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D4 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D5 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A1 = CLBLM_R_X5Y133_SLICE_X6Y133_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A2 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A5 = CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A6 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B1 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B2 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B4 = CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B6 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C2 = CLBLM_R_X5Y129_SLICE_X7Y129_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C3 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C5 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D5 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D5 = CLBLM_R_X5Y129_SLICE_X6Y129_D5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A1 = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A2 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A3 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A4 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A6 = CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_AX = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B1 = CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B2 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B3 = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B4 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B6 = CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B4 = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B5 = CLBLM_R_X7Y136_SLICE_X8Y136_CO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A3 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A4 = CLBLM_R_X3Y127_SLICE_X3Y127_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A5 = CLBLM_R_X7Y129_SLICE_X9Y129_C5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A1 = CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A2 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A3 = CLBLM_R_X5Y131_SLICE_X7Y131_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B1 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_AX = CLBLM_R_X5Y133_SLICE_X6Y133_DQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B2 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B1 = CLBLL_L_X4Y130_SLICE_X4Y130_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B2 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_DQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B4 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C2 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A1 = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A3 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A4 = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C3 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_DQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C5 = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D1 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D2 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D3 = CLBLM_L_X8Y126_SLICE_X11Y126_DQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D4 = CLBLL_L_X4Y127_SLICE_X4Y127_D5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D6 = CLBLM_R_X5Y132_SLICE_X6Y132_C5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A2 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A3 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A4 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_AX = CLBLM_L_X8Y126_SLICE_X11Y126_DQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B3 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C1 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C2 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C3 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C4 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C5 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C6 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D3 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D1 = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D2 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D3 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D6 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D3 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A1 = CLBLM_L_X8Y130_SLICE_X11Y130_D5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D4 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A4 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_CQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B1 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B2 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B3 = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B4 = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B5 = CLBLM_R_X11Y131_SLICE_X14Y131_CQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B6 = CLBLM_R_X11Y130_SLICE_X15Y130_A5Q;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C1 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C2 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C3 = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C4 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C6 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D3 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D4 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D5 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D6 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A2 = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A3 = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A4 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A6 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_AX = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B2 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B3 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B5 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B6 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C1 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C2 = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C4 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C5 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C6 = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D2 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D4 = CLBLL_L_X4Y129_SLICE_X4Y129_CQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D5 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A1 = CLBLL_L_X4Y127_SLICE_X4Y127_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A6 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_AX = CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B4 = CLBLM_L_X8Y127_SLICE_X11Y127_DQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B5 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B6 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A4 = CLBLM_R_X11Y127_SLICE_X14Y127_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A6 = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B1 = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B2 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B4 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B5 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A1 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C1 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C2 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C3 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C4 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C5 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C6 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A4 = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_C5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A6 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B1 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B5 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D1 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D4 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B6 = CLBLM_R_X5Y124_SLICE_X7Y124_B5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C2 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C4 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C6 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D2 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D4 = CLBLM_R_X5Y125_SLICE_X7Y125_C5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D5 = CLBLM_R_X7Y134_SLICE_X9Y134_B5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X13Y133_SLICE_X19Y133_AO5;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_AX = CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_BX = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = CLBLM_R_X11Y133_SLICE_X14Y133_DQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = CLBLM_R_X11Y131_SLICE_X14Y131_CQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = CLBLM_L_X8Y133_SLICE_X11Y133_CQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X4Y131_SLICE_X5Y131_C5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = CLBLM_R_X11Y131_SLICE_X14Y131_DQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A2 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_DQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A5 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B1 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B3 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B4 = CLBLM_L_X8Y134_SLICE_X11Y134_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B5 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C1 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C3 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C4 = CLBLM_L_X8Y130_SLICE_X10Y130_C5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D2 = CLBLM_R_X7Y128_SLICE_X9Y128_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D4 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D5 = CLBLM_L_X8Y129_SLICE_X10Y129_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A1 = CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A5 = CLBLM_L_X8Y130_SLICE_X11Y130_C5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A6 = CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B4 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B5 = CLBLM_L_X8Y128_SLICE_X10Y128_C5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B6 = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C2 = CLBLM_L_X8Y128_SLICE_X10Y128_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C3 = CLBLM_L_X10Y129_SLICE_X13Y129_C5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C5 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D1 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D2 = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D5 = CLBLM_R_X3Y127_SLICE_X2Y127_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A3 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A4 = CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A5 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B2 = CLBLM_L_X12Y127_SLICE_X16Y127_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B3 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B4 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B5 = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C2 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C3 = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C4 = CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C5 = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C6 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D2 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D4 = CLBLM_R_X11Y132_SLICE_X15Y132_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D5 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D6 = CLBLM_L_X10Y133_SLICE_X13Y133_D5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A1 = CLBLM_R_X7Y135_SLICE_X8Y135_DQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A2 = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A4 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A5 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B1 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B3 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B4 = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B5 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B6 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C2 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C4 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C5 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C6 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D1 = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D2 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D4 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D6 = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A1 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A2 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A3 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A5 = CLBLM_L_X10Y126_SLICE_X12Y126_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B1 = CLBLM_L_X8Y130_SLICE_X11Y130_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B2 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B6 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C1 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C2 = CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C3 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C5 = CLBLM_L_X10Y132_SLICE_X12Y132_DQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D1 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D3 = CLBLM_R_X3Y127_SLICE_X2Y127_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D4 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D5 = CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D6 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A1 = CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A2 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A3 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A4 = CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A5 = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B1 = CLBLM_L_X8Y133_SLICE_X11Y133_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B4 = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B5 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C1 = CLBLM_L_X8Y130_SLICE_X11Y130_C5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C5 = CLBLM_L_X12Y132_SLICE_X16Y132_DQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D3 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D5 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A1 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A3 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A4 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A6 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B1 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B2 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B4 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B5 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B6 = CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A1 = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A2 = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A4 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A5 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A6 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C1 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C2 = CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C3 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B1 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B2 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B5 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C3 = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C4 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C5 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C6 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D3 = CLBLM_L_X8Y134_SLICE_X10Y134_DQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A3 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A4 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D3 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D4 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D6 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A6 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B1 = CLBLM_R_X11Y132_SLICE_X15Y132_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B3 = CLBLM_R_X11Y133_SLICE_X14Y133_CQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B4 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A1 = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A2 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A4 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A6 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C1 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B1 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B2 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B3 = CLBLM_R_X5Y128_SLICE_X7Y128_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B4 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B6 = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C3 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D3 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D5 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D3 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D6 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C4 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = CLBLM_L_X8Y129_SLICE_X11Y129_CQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = CLBLL_L_X4Y132_SLICE_X4Y132_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = CLBLM_R_X5Y130_SLICE_X7Y130_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = CLBLM_R_X3Y131_SLICE_X3Y131_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = CLBLM_L_X8Y129_SLICE_X11Y129_CQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = CLBLM_L_X8Y131_SLICE_X11Y131_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = CLBLM_L_X8Y128_SLICE_X11Y128_C5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = CLBLM_R_X5Y125_SLICE_X7Y125_B5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B2 = CLBLM_L_X10Y129_SLICE_X13Y129_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B6 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A2 = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A4 = CLBLM_L_X10Y133_SLICE_X13Y133_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A6 = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B1 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B2 = CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B3 = CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B4 = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B6 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B4 = CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A1 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A2 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A3 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A4 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A6 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C2 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B1 = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B2 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B5 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_D5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C4 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C5 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C6 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D4 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A4 = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A5 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A6 = CLBLM_R_X11Y125_SLICE_X14Y125_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D3 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D4 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B1 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B2 = CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B4 = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B5 = CLBLM_R_X11Y134_SLICE_X14Y134_C5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A2 = CLBLM_R_X7Y128_SLICE_X8Y128_C5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A5 = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A6 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C2 = CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B1 = CLBLM_R_X5Y131_SLICE_X6Y131_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B3 = CLBLM_L_X10Y127_SLICE_X12Y127_B5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D1 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C1 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C3 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C4 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C5 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D3 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D4 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D1 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D3 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D4 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D5 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D6 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X11Y124_SLICE_X15Y124_B5Q;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X7Y131_SLICE_X9Y131_C5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D5 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = CLBLM_R_X7Y131_SLICE_X8Y131_D5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = CLBLM_R_X7Y135_SLICE_X8Y135_D5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = CLBLL_L_X4Y128_SLICE_X4Y128_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = CLBLM_L_X8Y129_SLICE_X10Y129_C5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_AX = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = CLBLM_R_X5Y131_SLICE_X6Y131_C5Q;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A2 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A4 = CLBLM_R_X3Y124_SLICE_X2Y124_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A5 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = CLBLM_L_X8Y131_SLICE_X11Y131_DQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = CLBLM_R_X7Y128_SLICE_X9Y128_CQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B2 = CLBLL_L_X2Y123_SLICE_X1Y123_BQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B4 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B5 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B6 = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C1 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C2 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C3 = CLBLL_L_X2Y123_SLICE_X1Y123_BQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C5 = CLBLM_R_X3Y124_SLICE_X2Y124_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C5 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C6 = CLBLM_L_X8Y129_SLICE_X10Y129_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A2 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A6 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B4 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B6 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = CLBLM_R_X7Y128_SLICE_X9Y128_C5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = CLBLM_L_X10Y125_SLICE_X12Y125_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A1 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A3 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A5 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = CLBLM_R_X7Y131_SLICE_X9Y131_C5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D6 = CLBLM_L_X8Y129_SLICE_X10Y129_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_AX = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B1 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B2 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B3 = CLBLM_R_X7Y133_SLICE_X8Y133_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C1 = CLBLM_R_X7Y133_SLICE_X8Y133_B5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C2 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C3 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = CLBLM_R_X5Y125_SLICE_X7Y125_B5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = CLBLM_L_X8Y128_SLICE_X11Y128_B5Q;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_L_X10Y125_SLICE_X13Y125_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = CLBLM_L_X8Y132_SLICE_X11Y132_B5Q;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = CLBLM_R_X7Y125_SLICE_X9Y125_B5Q;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A1 = CLBLM_L_X8Y133_SLICE_X11Y133_DQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A2 = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A3 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A5 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B1 = CLBLM_L_X8Y133_SLICE_X10Y133_D5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B2 = CLBLM_L_X8Y130_SLICE_X11Y130_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B4 = CLBLM_R_X5Y129_SLICE_X7Y129_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B5 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C1 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C3 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C4 = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C5 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D1 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D4 = CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D5 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A1 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A3 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_AX = CLBLM_R_X7Y125_SLICE_X9Y125_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B1 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B5 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_BX = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C1 = CLBLM_L_X8Y133_SLICE_X10Y133_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C2 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C3 = CLBLM_L_X8Y133_SLICE_X11Y133_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C4 = CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C5 = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C6 = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D2 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D3 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D4 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D6 = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A3 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A4 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A6 = CLBLM_R_X11Y125_SLICE_X14Y125_B5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B3 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B4 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A2 = CLBLM_L_X8Y125_SLICE_X11Y125_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A3 = CLBLM_R_X7Y128_SLICE_X9Y128_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A4 = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B2 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B3 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B5 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C1 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C2 = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C3 = CLBLM_R_X7Y126_SLICE_X9Y126_DQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C4 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D3 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A1 = CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A2 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A3 = CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A5 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D1 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D2 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D4 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D5 = CLBLM_R_X7Y124_SLICE_X9Y124_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B2 = CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B3 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B4 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B5 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B6 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B1 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A4 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A5 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A6 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C1 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C2 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C3 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B5 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B6 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D2 = CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C2 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C4 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C5 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D3 = CLBLM_L_X10Y126_SLICE_X12Y126_DQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D6 = CLBLM_R_X11Y125_SLICE_X14Y125_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D1 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D2 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D3 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D4 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D5 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = CLBLM_R_X11Y132_SLICE_X15Y132_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = CLBLM_R_X5Y132_SLICE_X6Y132_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = CLBLM_R_X7Y133_SLICE_X9Y133_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = CLBLM_L_X8Y133_SLICE_X11Y133_CQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = CLBLM_L_X8Y135_SLICE_X11Y135_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = CLBLM_R_X5Y131_SLICE_X7Y131_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = CLBLM_L_X8Y133_SLICE_X11Y133_DQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = CLBLM_R_X7Y133_SLICE_X9Y133_DQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = CLBLM_L_X8Y132_SLICE_X11Y132_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = CLBLM_L_X8Y134_SLICE_X10Y134_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = CLBLM_L_X8Y130_SLICE_X10Y130_DQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A1 = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A2 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A3 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A6 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B1 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B3 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B5 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B6 = CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C1 = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C4 = CLBLL_L_X4Y128_SLICE_X5Y128_D5Q;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C5 = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A1 = CLBLM_R_X11Y126_SLICE_X15Y126_B5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A2 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A3 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D3 = CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D4 = CLBLM_R_X7Y127_SLICE_X9Y127_DQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D6 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A1 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A2 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A4 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A5 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_AX = CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B1 = CLBLM_R_X5Y128_SLICE_X7Y128_C5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B3 = CLBLM_L_X8Y129_SLICE_X10Y129_DQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B5 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_BX = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C1 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C3 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C5 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C6 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D2 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D5 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D6 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A2 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A4 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A6 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B1 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B2 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B4 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B5 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B6 = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C2 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C3 = CLBLM_L_X8Y132_SLICE_X11Y132_DQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C5 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D2 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D3 = CLBLM_L_X8Y134_SLICE_X11Y134_DQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D4 = CLBLM_L_X8Y130_SLICE_X11Y130_DQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D5 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A1 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A2 = CLBLM_L_X8Y134_SLICE_X10Y134_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A3 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_D5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_AX = CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B1 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B2 = CLBLM_L_X8Y134_SLICE_X10Y134_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B5 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B6 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C4 = CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C5 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D1 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D2 = CLBLM_L_X8Y134_SLICE_X10Y134_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D4 = CLBLM_L_X8Y134_SLICE_X11Y134_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A1 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A2 = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A4 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A6 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B1 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B2 = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B4 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B5 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C1 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C2 = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C4 = CLBLM_R_X11Y128_SLICE_X14Y128_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C5 = CLBLM_R_X3Y129_SLICE_X3Y129_DQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D2 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D4 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D5 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A1 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A3 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A4 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A6 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y194_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B1 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B2 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B4 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B6 = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign LIOB33_X0Y193_IOB_X0Y193_O = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C1 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C2 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C5 = CLBLL_L_X4Y128_SLICE_X5Y128_CQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D2 = CLBLL_L_X4Y127_SLICE_X5Y127_DQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D4 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D6 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C4 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B4 = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B6 = CLBLM_R_X13Y133_SLICE_X18Y133_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A1 = CLBLM_L_X8Y134_SLICE_X11Y134_DQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A3 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A5 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A6 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B1 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B2 = CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B4 = CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B6 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C2 = CLBLM_L_X10Y125_SLICE_X13Y125_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C4 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C5 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D1 = CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D2 = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D3 = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D4 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D5 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C6 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A2 = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A3 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A4 = CLBLM_R_X7Y135_SLICE_X9Y135_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A5 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_AX = CLBLM_L_X8Y129_SLICE_X10Y129_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B2 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C1 = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C2 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C3 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C5 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D1 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D2 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D3 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D5 = CLBLM_L_X10Y135_SLICE_X13Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D6 = CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A6 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D5 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_AX = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = CLBLL_L_X4Y126_SLICE_X5Y126_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_C5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = CLBLM_R_X7Y131_SLICE_X9Y131_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_B5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = CLBLL_L_X4Y128_SLICE_X4Y128_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_DQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = CLBLL_L_X4Y128_SLICE_X5Y128_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C4 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C5 = CLBLM_L_X8Y132_SLICE_X11Y132_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C6 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = CLBLM_L_X8Y125_SLICE_X10Y125_C5Q;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A3 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = CLBLM_R_X5Y131_SLICE_X6Y131_CQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A5 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B5 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C5 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = CLBLM_L_X12Y132_SLICE_X16Y132_D5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A1 = CLBLM_L_X10Y126_SLICE_X12Y126_DQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A3 = CLBLM_R_X11Y125_SLICE_X14Y125_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A4 = CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B1 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B3 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B6 = CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C5 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D5 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A1 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A2 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A4 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A5 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B2 = CLBLM_L_X8Y125_SLICE_X10Y125_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B3 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B4 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B5 = CLBLM_R_X11Y133_SLICE_X14Y133_CQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C1 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C2 = CLBLM_R_X5Y128_SLICE_X7Y128_CQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C3 = CLBLL_L_X2Y123_SLICE_X1Y123_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C5 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D1 = CLBLM_R_X3Y127_SLICE_X3Y127_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D2 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D3 = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A4 = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A6 = CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B1 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B2 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B3 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B4 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B5 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C3 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C5 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C6 = CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D6 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = CLBLM_R_X5Y126_SLICE_X6Y126_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_AX = CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = CLBLM_R_X7Y130_SLICE_X9Y130_DQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = CLBLM_R_X5Y131_SLICE_X7Y131_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = CLBLM_L_X8Y134_SLICE_X10Y134_CQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = CLBLM_L_X8Y129_SLICE_X10Y129_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = CLBLM_L_X10Y133_SLICE_X12Y133_DQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = CLBLM_R_X5Y132_SLICE_X6Y132_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C2 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = CLBLM_R_X7Y131_SLICE_X9Y131_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = CLBLM_L_X8Y128_SLICE_X11Y128_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = CLBLM_R_X7Y133_SLICE_X9Y133_DQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = CLBLM_L_X8Y127_SLICE_X10Y127_DQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = CLBLM_R_X11Y124_SLICE_X15Y124_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = CLBLM_R_X7Y133_SLICE_X9Y133_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_AX = CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = CLBLM_R_X3Y130_SLICE_X2Y130_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = CLBLM_L_X8Y133_SLICE_X10Y133_DQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D4 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C5 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C4 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign LIOB33_X0Y195_IOB_X0Y196_O = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign LIOB33_X0Y195_IOB_X0Y195_O = CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A2 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A6 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A2 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A3 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A6 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B1 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B2 = CLBLM_R_X7Y131_SLICE_X8Y131_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B3 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B5 = CLBLM_R_X7Y126_SLICE_X9Y126_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D2 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C2 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C3 = CLBLM_R_X7Y130_SLICE_X9Y130_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C5 = CLBLM_L_X8Y133_SLICE_X10Y133_DQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D2 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D3 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D4 = CLBLM_L_X8Y134_SLICE_X10Y134_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D5 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A1 = CLBLM_R_X7Y133_SLICE_X8Y133_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A3 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A4 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A5 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B1 = CLBLM_L_X8Y133_SLICE_X10Y133_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B3 = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B5 = CLBLM_R_X7Y132_SLICE_X8Y132_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D5 = CLBLM_L_X8Y130_SLICE_X10Y130_D5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B4 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C1 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C3 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C6 = CLBLM_R_X5Y133_SLICE_X7Y133_D5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B6 = CLBLM_L_X8Y128_SLICE_X11Y128_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D2 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D5 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X4Y127_SLICE_X5Y127_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C5 = CLBLM_R_X7Y126_SLICE_X8Y126_C5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B5 = CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B6 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = CLBLM_R_X5Y128_SLICE_X7Y128_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A1 = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A2 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A3 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A4 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B3 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B4 = CLBLM_R_X11Y128_SLICE_X14Y128_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B5 = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A2 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A3 = CLBLL_L_X4Y128_SLICE_X5Y128_DQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C2 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C3 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B1 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B2 = CLBLL_L_X4Y124_SLICE_X5Y124_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B5 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D1 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C1 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C2 = CLBLM_L_X8Y130_SLICE_X10Y130_B5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C3 = CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C5 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C6 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D4 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A1 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A3 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A4 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D1 = CLBLL_L_X4Y124_SLICE_X5Y124_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D2 = CLBLM_L_X8Y128_SLICE_X10Y128_DQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D3 = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D4 = CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D6 = CLBLM_R_X3Y127_SLICE_X2Y127_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A6 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B1 = CLBLM_R_X7Y129_SLICE_X9Y129_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B2 = CLBLM_R_X7Y131_SLICE_X8Y131_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B4 = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A1 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A2 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A4 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C1 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C2 = CLBLM_R_X11Y133_SLICE_X14Y133_DQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B1 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B2 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B4 = CLBLM_R_X5Y127_SLICE_X6Y127_C5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D2 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D3 = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C5 = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D4 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D5 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D6 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C5 = CLBLM_R_X11Y134_SLICE_X14Y134_B5Q;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = CLBLL_L_X4Y127_SLICE_X4Y127_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C6 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = CLBLM_R_X3Y128_SLICE_X3Y128_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A2 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A3 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A4 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A5 = CLBLM_R_X7Y134_SLICE_X9Y134_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A6 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_AX = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B2 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B3 = CLBLM_L_X8Y130_SLICE_X11Y130_DQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B4 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B5 = CLBLM_R_X7Y133_SLICE_X9Y133_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B6 = CLBLM_L_X8Y131_SLICE_X11Y131_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_BX = CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A1 = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A3 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A4 = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A5 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C2 = CLBLM_R_X7Y135_SLICE_X9Y135_CQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C4 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B1 = CLBLL_L_X4Y128_SLICE_X5Y128_DQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B2 = CLBLM_R_X7Y128_SLICE_X8Y128_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B4 = CLBLM_R_X5Y127_SLICE_X6Y127_D5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C3 = CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C4 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D3 = CLBLM_R_X11Y125_SLICE_X14Y125_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D4 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A1 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A2 = CLBLM_R_X7Y135_SLICE_X8Y135_DQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A3 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A5 = CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D2 = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D4 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A6 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B3 = CLBLM_R_X7Y132_SLICE_X8Y132_C5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B4 = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A1 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A2 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A4 = CLBLM_R_X5Y128_SLICE_X6Y128_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C1 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C2 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_B5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B2 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B5 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B6 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D1 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C2 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C4 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C5 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C6 = CLBLL_L_X4Y127_SLICE_X5Y127_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D3 = CLBLM_L_X8Y130_SLICE_X10Y130_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D1 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D2 = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D4 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D5 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D6 = 1'b1;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A1 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A2 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A5 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A6 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B1 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B3 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B4 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B6 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C1 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C2 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = CLBLL_L_X4Y128_SLICE_X4Y128_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_D5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D3 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D4 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A1 = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A2 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A3 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A5 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_DQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = CLBLM_L_X8Y134_SLICE_X11Y134_D5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A6 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B1 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B4 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B2 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = CLBLL_L_X4Y127_SLICE_X4Y127_B5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = CLBLL_L_X4Y126_SLICE_X5Y126_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C1 = CLBLM_L_X8Y135_SLICE_X11Y135_C5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = CLBLM_R_X7Y128_SLICE_X9Y128_DQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_D5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D1 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D2 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = CLBLM_R_X7Y130_SLICE_X9Y130_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D5 = CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D6 = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = CLBLL_L_X4Y128_SLICE_X5Y128_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D5 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A2 = CLBLM_R_X7Y136_SLICE_X9Y136_DO5;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A6 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = CLBLM_R_X5Y133_SLICE_X6Y133_C5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = CLBLM_R_X5Y129_SLICE_X7Y129_CQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = CLBLM_L_X8Y129_SLICE_X11Y129_DQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A2 = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A3 = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A4 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A5 = CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = CLBLM_R_X7Y128_SLICE_X9Y128_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B3 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = CLBLL_L_X4Y127_SLICE_X4Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = CLBLM_L_X8Y128_SLICE_X11Y128_C5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = CLBLL_L_X4Y127_SLICE_X5Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = CLBLL_L_X4Y126_SLICE_X5Y126_A5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = CLBLM_L_X8Y134_SLICE_X11Y134_C5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B6 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_DQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A4 = CLBLM_R_X7Y127_SLICE_X9Y127_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B1 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B2 = CLBLM_R_X5Y125_SLICE_X7Y125_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B5 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C1 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C2 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C5 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D2 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D3 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A3 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A4 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A5 = CLBLM_R_X11Y133_SLICE_X14Y133_D5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B3 = CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B5 = CLBLM_R_X3Y127_SLICE_X3Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B6 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C1 = CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C4 = CLBLM_R_X7Y128_SLICE_X8Y128_D5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C5 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D1 = CLBLL_L_X4Y129_SLICE_X5Y129_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D4 = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C4 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C5 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
endmodule
