module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD
  );
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BQ;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CLK;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CLK;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CQ;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CLK;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AQ;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BQ;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CLK;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CQ;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AQ;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CLK;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CQ;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AQ;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CLK;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CE;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5Q;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CLK;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5Q;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CLK;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CLK;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CLK;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CLK;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CLK;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5Q;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CLK;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CLK;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CLK;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CLK;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CLK;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CLK;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.Q(CLBLL_L_X2Y108_SLICE_X1Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.Q(CLBLL_L_X2Y108_SLICE_X1Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff888888ff882888)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(CLBLL_L_X2Y109_SLICE_X1Y109_DO6),
.I1(CLBLL_L_X2Y108_SLICE_X1Y108_BQ),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_AQ),
.I3(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heca0eca0ce0ace0a)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(CLBLL_L_X2Y109_SLICE_X1Y109_DO6),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaababaaa00ba20)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_CQ),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0300aaaa03ff)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_CQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050404050004040)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_CQ),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f0070778f88)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I4(CLBLL_L_X2Y109_SLICE_X1Y109_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y109_SLICE_X1Y109_AO6),
.Q(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y109_SLICE_X1Y109_BO6),
.Q(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y109_SLICE_X1Y109_CO6),
.Q(CLBLL_L_X2Y109_SLICE_X1Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f50f0a0f0a)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3caa00be3caa00)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_CQ),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y109_SLICE_X1Y109_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0e4a0b4a0b4)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_AQ),
.I3(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.I4(1'b1),
.I5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haabe00503f3fffff)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I3(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.I4(CLBLL_L_X2Y109_SLICE_X1Y109_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.Q(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555500000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0f5f0faa00aa00)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff00c6cc0000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_CQ),
.I1(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I4(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55551111f5fff1f3)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff3fffffffb)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I1(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.I5(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fc00a8ffffaafe)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_CO6),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_DO6),
.I3(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_BQ),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8ccc8ccc8cc3233)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_CO6),
.I1(CLBLL_L_X2Y108_SLICE_X1Y108_BQ),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_DO6),
.I3(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I4(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f06636cc3c)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.I1(CLBLL_L_X2Y108_SLICE_X1Y108_BQ),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.Q(CLBLL_L_X2Y111_SLICE_X0Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.Q(CLBLL_L_X2Y111_SLICE_X0Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.Q(CLBLL_L_X2Y111_SLICE_X0Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaffafafaf9)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_CQ),
.I2(CLBLL_L_X2Y111_SLICE_X0Y111_BQ),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_AQ),
.I4(CLBLL_L_X2Y111_SLICE_X0Y111_AQ),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_CQ),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffecececffa0a0a0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_CQ),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefaeeaafcf0cc00)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_BQ),
.I2(CLBLL_L_X2Y111_SLICE_X0Y111_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X2Y111_SLICE_X0Y111_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AQ),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff0f0f0f0)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y111_SLICE_X0Y111_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aa8aa080)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_CQ),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bdeffffffff7bde)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(CLBLL_L_X2Y111_SLICE_X0Y111_AQ),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_AQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I5(CLBLL_L_X2Y111_SLICE_X0Y111_CQ),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccf33303330)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.Q(CLBLL_L_X2Y112_SLICE_X0Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y112_SLICE_X0Y112_BO6),
.Q(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.Q(CLBLL_L_X2Y112_SLICE_X0Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d050d05020a020a)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefceeccfaf0aa00)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_CQ),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefaeeaafcf0cc00)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff888f888f888)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.Q(CLBLL_L_X2Y112_SLICE_X1Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfc0cfc0c)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h777c7478777c7478)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_A5Q),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404c2c205050101)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101a0a000004444)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444088444e4088)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_CQ),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_A5Q),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf098f00023232323)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_A5Q),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa1ff0000a10000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_A5Q),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfefdfeffdfefdfe)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3100000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc07cc08cc0fcc00)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff410050ff410050)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55fffdff55fff5ff)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000066004400)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff10ffc0001000c0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_CQ),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_A5Q),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb100b177777777)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000330000001300)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcfaf0cecc0a00)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_BQ),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0d0d00000d0d)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccca04400005555)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf90cf000bbffbbff)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_A5Q),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_A5Q),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaea4040bbbb0000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f000a0a0c0c)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_A5Q),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30b03030ff55ffff)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088f020f088)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa000a0ff0200a0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000550000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haac3aa00aac3aa00)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa330f33aa330f33)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77f333f3fff333f3)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff2f20efe0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff62ffaa00400000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f8fff8f0f0fff0f)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b888b88b888b8)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hef00ff00ff00ff00)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7f00000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aac3aa00aac3)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffffffffff)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfff5fffffffff)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7fff7fff7ff)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff300030ff030030)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfff8fffcfffcf)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033333233)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_BQ),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceedcdc00221010)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_BQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_DQ),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeffcccccccc)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0aca3a0a0a6a3)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c0009ff0c0009)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0082a0ff00a0a0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_DO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fdfff0f0f2f0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_CQ),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff00ffccffa0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f888888888f8f8)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00000c000a0a)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_CQ),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.Q(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaffafafaf5)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_CQ),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5151404011110000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0cc00f0f0aaaa)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_DQ),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_AQ),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff022f000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_CQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcccccccfcccdcc)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_DO6),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.I2(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff03ff0fff03ff0b)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_DO6),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_BO6),
.I2(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7070007008080f08)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_CQ),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_AQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88ff88888fff8f8f)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccdcdcccc)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff040000ff04)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb4bbbaaaa5aaa)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88cc0000c8c80000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.Q(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.Q(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.Q(CLBLM_R_X3Y111_SLICE_X2Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0c0f0f0a0c0a)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8888ff88888888)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_CQ),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404f104f104)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_BQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5014ff3fff3f)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaa200008880)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_CQ),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_BQ),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04fa00fa00fa00)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c8c8c8c0c8c8c8)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0aa00eecceecc)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.Q(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.Q(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.Q(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.Q(CLBLM_R_X3Y112_SLICE_X2Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2c0c0e2e2c0c0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaeaffff0040)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_DQ),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaafaffaaeaea)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_DQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff005a5a)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_A5Q),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccecccccccccc8)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_AQ),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef4041111bbbb)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_A5Q),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4f0f044440000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_BQ),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05055555ea40ea40)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff90c00000c0c0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaffaafafabbaa)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_DQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hecec0220ecec0220)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000eeccaa00)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.I2(1'b1),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcc00ffffcc40)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff04a4000004a4)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_A5Q),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000505ff000505)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa003caaaa003c)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha6aca6aca0a0a0a0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_CQ),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I4(1'b1),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001230ff001230)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeaaaffaaaaaaff)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_CQ),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5fffff5f577ff)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_A5Q),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ffffff75ffffff)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_CQ),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_A5Q),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h40ff0000bf00bf00)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_A5Q),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_A5Q),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00bfbfffffbfbf)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f00aaaa0008)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f04444f0f00014)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff404100004041)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_CQ),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc50cc50cc50cc41)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.Q(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff70ffff)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00020202ffffffff)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8cff0cffccffcc)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00e105050505)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_CO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff77ff00ff)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000c0c0303)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808f808f202f202)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000050055005)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdf)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005000700050005)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_CQ),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_CO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777700800000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa5000000a500)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc88888888d8d8)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaaee00000044)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff414100004141)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0cc28cca0cc28)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_R_X3Y113_SLICE_X3Y113_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_AMUX = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_BMUX = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_AMUX = CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_DMUX = CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_AMUX = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_CMUX = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_AMUX = CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_AMUX = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_DMUX = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D = CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_AMUX = CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_BMUX = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_AMUX = CLBLL_L_X4Y108_SLICE_X4Y108_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_BMUX = CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_DMUX = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_AMUX = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_AMUX = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_AMUX = CLBLL_L_X4Y110_SLICE_X5Y110_A5Q;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_BMUX = CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_CMUX = CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_DMUX = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_CMUX = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_DMUX = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_BMUX = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_DMUX = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_AMUX = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_BMUX = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_DMUX = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AMUX = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_BMUX = CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_AMUX = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_DMUX = CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_A5Q;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_BMUX = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_CMUX = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_DMUX = CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_AMUX = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_AMUX = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_DMUX = CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_AMUX = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_BMUX = CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = CLBLL_L_X2Y111_SLICE_X0Y111_BQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = CLBLL_L_X2Y111_SLICE_X0Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = CLBLL_L_X2Y111_SLICE_X0Y111_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = CLBLL_L_X2Y111_SLICE_X0Y111_BQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = CLBLL_L_X2Y111_SLICE_X0Y111_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = CLBLL_L_X2Y111_SLICE_X0Y111_BQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = CLBLL_L_X2Y112_SLICE_X0Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = CLBLL_L_X2Y111_SLICE_X0Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = CLBLM_R_X3Y111_SLICE_X2Y111_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = CLBLL_L_X2Y111_SLICE_X0Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = CLBLL_L_X2Y112_SLICE_X0Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = CLBLL_L_X2Y111_SLICE_X0Y111_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = CLBLL_L_X2Y112_SLICE_X0Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = CLBLL_L_X4Y110_SLICE_X5Y110_A5Q;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = CLBLL_L_X2Y112_SLICE_X0Y112_AQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = CLBLL_L_X2Y112_SLICE_X0Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = CLBLM_R_X3Y112_SLICE_X2Y112_DQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = CLBLM_R_X3Y109_SLICE_X2Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = CLBLM_R_X3Y109_SLICE_X2Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = CLBLM_R_X3Y109_SLICE_X2Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = CLBLL_L_X4Y108_SLICE_X4Y108_CQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = CLBLM_R_X3Y109_SLICE_X3Y109_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = CLBLL_L_X2Y111_SLICE_X0Y111_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = CLBLL_L_X2Y112_SLICE_X0Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = CLBLM_R_X3Y111_SLICE_X2Y111_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = CLBLL_L_X2Y112_SLICE_X0Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = CLBLM_R_X3Y112_SLICE_X3Y112_A5Q;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = CLBLL_L_X2Y112_SLICE_X1Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = CLBLL_L_X2Y112_SLICE_X1Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = CLBLL_L_X4Y109_SLICE_X5Y109_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_A5Q;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = CLBLM_R_X3Y112_SLICE_X2Y112_DQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = CLBLM_R_X3Y112_SLICE_X2Y112_DQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = CLBLL_L_X2Y112_SLICE_X0Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_AX = CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = CLBLL_L_X4Y110_SLICE_X5Y110_A5Q;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLL_L_X4Y109_SLICE_X5Y109_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLL_L_X4Y110_SLICE_X5Y110_A5Q;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLL_L_X4Y108_SLICE_X4Y108_A5Q;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = CLBLM_R_X3Y112_SLICE_X2Y112_DQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = CLBLL_L_X4Y109_SLICE_X5Y109_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_CE = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = CLBLM_R_X3Y111_SLICE_X3Y111_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = CLBLL_L_X4Y108_SLICE_X4Y108_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_AX = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = CLBLL_L_X4Y108_SLICE_X4Y108_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = CLBLL_L_X4Y108_SLICE_X4Y108_CQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AX = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = CLBLL_L_X4Y108_SLICE_X4Y108_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = CLBLM_R_X3Y109_SLICE_X2Y109_DQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = CLBLL_L_X4Y109_SLICE_X5Y109_CQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = CLBLL_L_X4Y110_SLICE_X5Y110_A5Q;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = CLBLL_L_X2Y108_SLICE_X1Y108_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = CLBLL_L_X2Y109_SLICE_X1Y109_CQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = CLBLL_L_X2Y108_SLICE_X1Y108_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = CLBLL_L_X2Y112_SLICE_X0Y112_CQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = CLBLL_L_X2Y112_SLICE_X0Y112_CQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = CLBLL_L_X2Y112_SLICE_X0Y112_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = CLBLL_L_X2Y109_SLICE_X1Y109_CQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_AX = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = CLBLL_L_X4Y110_SLICE_X5Y110_A5Q;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = CLBLL_L_X4Y108_SLICE_X4Y108_A5Q;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = CLBLL_L_X2Y109_SLICE_X1Y109_CQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = CLBLL_L_X2Y108_SLICE_X1Y108_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = CLBLL_L_X2Y109_SLICE_X1Y109_CQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = CLBLM_R_X3Y111_SLICE_X2Y111_CQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = CLBLM_R_X3Y111_SLICE_X2Y111_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = CLBLL_L_X2Y108_SLICE_X1Y108_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = CLBLL_L_X2Y108_SLICE_X1Y108_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = CLBLL_L_X2Y108_SLICE_X1Y108_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = CLBLM_R_X3Y112_SLICE_X2Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = CLBLL_L_X2Y111_SLICE_X0Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = CLBLL_L_X2Y112_SLICE_X0Y112_AQ;
endmodule
