module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CLK;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5Q;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CLK;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AMUX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AMUX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_BO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_BO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_DO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AMUX;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CLK;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CLK;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5Q;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5Q;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CLK;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B5Q;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5Q;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CE;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_SR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5Q;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5Q;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DMUX;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5Q;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CE;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_SR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CLK;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CLK;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_DO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CLK;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_DO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CLK;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_AO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_AO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_BO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_BO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CLK;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_DO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_DO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AMUX;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_BO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_BO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_CO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_CO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_DO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C5Q;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CLK;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D5Q;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CLK;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CE;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_SR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CMUX;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AMUX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CE;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_SR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CLK;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5Q;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CLK;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5Q;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CLK;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5Q;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5Q;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C5Q;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5Q;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D5Q;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AMUX;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AMUX;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CLK;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CLK;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A5Q;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DMUX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CE;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_SR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AMUX;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_BO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_BO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CLK;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_DO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_DO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_BO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_BO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_CO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_CO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_DO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_DO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CLK;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AMUX;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_DO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CLK;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DMUX;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_BO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_DO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CLK;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CMUX;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_DO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_DO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BMUX;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CMUX;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_XOR;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A1;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A2;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A3;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A4;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_AMUX;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_AO5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_AO6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A_CY;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_A_XOR;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B1;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B2;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B3;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B4;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_BO5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_BO6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B_CY;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_B_XOR;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C1;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C2;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C3;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C4;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_CO5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_CO6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C_CY;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_C_XOR;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D1;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D2;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D3;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D4;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_DO5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_DO6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D_CY;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X42Y141_D_XOR;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A1;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A2;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A3;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A4;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_AO5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_AO6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A_CY;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_A_XOR;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B1;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B2;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B3;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B4;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_BO5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_BO6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B_CY;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_B_XOR;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C1;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C2;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C3;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C4;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_CO5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_CO6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C_CY;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_C_XOR;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D1;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D2;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D3;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D4;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_DO5;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_DO6;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D_CY;
  wire [0:0] CLBLM_R_X29Y141_SLICE_X43Y141_D_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_AO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_A_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_BO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_BO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_B_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_CO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_CO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_C_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_DO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_DO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X56Y120_D_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_AO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_AO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_A_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_BO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_BO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_B_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_CO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_CO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_C_XOR;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D1;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D2;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D3;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D4;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_DO5;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_DO6;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D_CY;
  wire [0:0] CLBLM_R_X37Y120_SLICE_X57Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5Q;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CLK;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CLK;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CLK;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CLK;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5Q;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5Q;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CLK;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CLK;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CLK;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CLK;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5Q;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CLK;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CLK;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5Q;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5Q;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AMUX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CLK;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5Q;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CLK;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5Q;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CLK;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5Q;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D5Q;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffdfffffffdfd)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffdfffffdfd)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc55550000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_CLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfbfffffffaf)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeffffffeeffff)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcddfd00f055f5)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc80cc80cc80)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_BO6),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_C5Q),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.Q(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaaafffcffff)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88bb88b888b8)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.Q(CLBLL_L_X2Y119_SLICE_X1Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.Q(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0cfcfffff)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_CQ),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_A5Q),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccffcc00cc00)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccdfcfddcc)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I1(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_BQ),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8c8c8c8c8cff8c8c)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7f5fffff3f0)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_BO6),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff0cffffffae)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I3(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff3f0fbfa)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffff7fffffff)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffaaee)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000008)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.I3(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_CO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003200000010)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I3(CLBLM_R_X29Y141_SLICE_X42Y141_AO6),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(LIOB33_X0Y61_IOB_X0Y61_I),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0fafffff0fa)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_BQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_CO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffffddffffff)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffffffff7ffff)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffffffffffef)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffffffeff)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000330050507350)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_CLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I2(LIOB33_X0Y57_IOB_X0Y57_I),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I4(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I5(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(LIOB33_X0Y53_IOB_X0Y54_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfffffdffffff)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_DLUT (
.I0(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_DO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_CLUT (
.I0(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_CO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000223000)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLM_R_X29Y141_SLICE_X42Y141_AO6),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_BO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddffffffffbbbb)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000220000002200)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_BO6),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_DO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdf)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_CLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_BO6),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_AO6),
.I5(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_CO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d0c5d0cffff5d0c)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I1(LIOB33_X0Y67_IOB_X0Y68_I),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_BO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c00cf00f05050)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_ALUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_AO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffff)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000303000001030)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLL_L_X2Y124_SLICE_X1Y124_AO6),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_BO6),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_CO6),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0008008dfffffff)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_ALUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfabafaba50105010)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccaaaa0c0c)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_B5Q),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaae000400f000f0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff770077ff700070)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880077777777)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a0afa0ac)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_DO6),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0cfccccc)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddd8d8d8d8)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaff000030303030)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_C5Q),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_A5Q),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haacfaa00aa03aa00)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f088882222)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaccaaccf0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffddddffffffff)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfffffffffff)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_DQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000570000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_C5Q),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2f3c0c0d1c0c0c0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_DQ),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_CO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaacccc00ff)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000006c006c)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00005550)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f5fff5f3300ff00)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdffffff)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa00c0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heecceecceac0eac0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffff0000ffff)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0f5a0f5a0a0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_A5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f101f404f404)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_B5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff120012ff120012)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0c0c0c0c0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaf0005afaa0500)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f808f000f000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_CO6),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc50ccffccf0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_C5Q),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc8c00cccc8c8c)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_DO6),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccf0ccf0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y127_IOB_X1Y127_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf8fff00d080f00)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_A5Q),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcdc3010ffdf3313)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_A5Q),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I5(LIOB33_X0Y53_IOB_X0Y53_I),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_BO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_DO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044aabb0011)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeaeae54540404)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I3(1'b1),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ff00fcf0cc00)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0f0affaa)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc800c8fffa00fa)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaf0aaf0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aa00aaf0aa00)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fa50fa50)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_C5Q),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffffc)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.I2(CLBLM_R_X5Y120_SLICE_X7Y120_B5Q),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ccaaccaa)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_C5Q),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I4(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf3aaffaac0aa00)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcf0fcf00cc00cc)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_CQ),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7f3f5f0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d00080000000000)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_DO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefafefacc00cc00)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_B5Q),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000c0a0a000c)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03030a0000000a00)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I2(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aac0aaffaacc)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00b8b8ff00b8b8)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffae)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_AO6),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_DO6),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_CO6),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_CLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.I3(CLBLL_L_X2Y124_SLICE_X1Y124_CO6),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f444f00004444)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_ALUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I4(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000000)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010000000)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaafaeefe)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfff0ff5a)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50ff505050ff5050)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_DLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fff5ff00fff0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_CLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfbbbfbaafaaafa)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_BLUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_DO6),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y55_IOB_X0Y55_I),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_ALUT (
.I0(CLBLL_L_X4Y123_SLICE_X5Y123_CO6),
.I1(CLBLL_L_X2Y124_SLICE_X1Y124_CO6),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h444400004f440f00)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I3(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaeffaeae)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_CLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_AO6),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I5(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000000000000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300030023222322)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I3(LIOB33_X0Y69_IOB_X0Y70_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa000c)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_DQ),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdc)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_BLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I3(CLBLL_L_X4Y123_SLICE_X4Y123_DO6),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_AO6),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_CO6),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202020202ff0202)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f20002)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_DLUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_B5Q),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeefffe)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_CLUT (
.I0(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I1(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_DO6),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002222f000f222)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_DQ),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I4(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h555d000c000c000c)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_ALUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_CQ),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I4(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfefcfefcceeccee)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_DLUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_BO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_A5Q),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_BLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_DO6),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_DO6),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_BO6),
.I5(CLBLL_L_X2Y124_SLICE_X1Y124_CO6),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfdffffff)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b0a3b0a3b0a3b0a)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdc)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_CLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_CO6),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BO6),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_CO6),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_BO6),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f200000002)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_BLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa00fa00)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000aac0c0c0ea)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_CLUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_A5Q),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3ffffff3fffff)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdefc1230fcfc3030)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcdc50505050)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_A5Q),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880088008800)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h400000004000c000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0aff08000a0008)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_A5Q),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcdddcd11011101)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c000f03000c030f)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_CQ),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_B5Q),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0a0a0a0a0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88b88800000f0f)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_DQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc50cc50cc55cc55)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_DO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc00fc00)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_A5Q),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00cc00)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y114_SLICE_X11Y114_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f011f055f011)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00ff00cc)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ff00c0c0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_DQ),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33003000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_BO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ff33ff3cffccffc)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0c00ffff0c)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_DO6),
.I3(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_B5Q),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f404f404)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a0f0a00f5f0f5f)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_DLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff03570357)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff11f111)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f033f000f000)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000900900009009)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_DLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_C5Q),
.I4(CLBLM_L_X8Y114_SLICE_X11Y114_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2100000000210000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_CLUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_B5Q),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3caaaa3f3caaaa)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_DO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff33fc30)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_CQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_DQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_DO6),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550055fffffff3)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccff500050)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I1(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_A5Q),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0c0c0eeee2222)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccde0012cdec0120)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_DLUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CQ),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.I5(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc0c0cc88cc88)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8d8d8d88888888)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54fe54aa00)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaa0ccccfff0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_DQ),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_DQ),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088ccffcc00)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000e0eff000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44ee44fa50)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e0d0e0e0e0e0e0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a020aaaaa0a0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee0000ff00f0f0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88dd88ddd8d8)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a020aaaa)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cf000fc0cf000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaf5005fbae5104)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.I3(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005555ff005050)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_ALUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_BO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_CO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f070f0f80008)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0aca0a0a0aca0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hababaeae01010404)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaeaffff5040)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_CO6),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_B5Q),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_BO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_CO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_DO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccf0ccaacca0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f808f000f808)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefaea55445040)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafffa00005550)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfeccce03030303)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff004444ccccf0f0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000bebe1414)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.I3(1'b1),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888dd8888dd88)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_CO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_DO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccff00c0c0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_DQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_CO6),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cc0cac0ca)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000bbee1144)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50aa00fa50)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_C5Q),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffffffff)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffff)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_CLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000200000)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff300030ff300030)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_CO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000101000001010)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_DLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00f000c0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0c0eeee2222)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_CO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_DO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcecccccfcec)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca0a0a0a0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_CLUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5e4a0a0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeaffeaaaeaaaea)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_CO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_DQ),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0fff000)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc55cc55cc00)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecc3200fa00fa00)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_BO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_CO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacafa0afa0a)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_DLUT (
.I0(RIOB33_X105Y143_IOB_X1Y144_I),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fafa0a0a)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5a0ccccf5a0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_ALUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_DLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc03fc738f00ff708)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_CLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff1f0f11001100)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_CO6),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_CO6),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa300c0330)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_ALUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_DQ),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_DO5),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_DO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dd88dd88)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbe00bec0c0c0c0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa03aa0caa0caa0c)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3fffaaaaffff)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_D5Q),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_CO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_BO5),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010ffff1010ffff)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_DLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fd000f000c00)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_CLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h08080000f5f00500)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_CQ),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd8888d8ddd888)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I5(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333332300000050)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f50505f0f00000)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_DQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccaaf0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h26f62727b505b5b5)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d888d888d888d88)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05511f0f00044)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000075207520)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fc30fc30)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0bbbbbbbb)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac0cc00cc00cc)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_DQ),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3fffffa000a000)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y141_I),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y139_IOB_X1Y140_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50000000ccccc6cc)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdddd0f0f0f87)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f0fffff8000ffff)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccedcc00002100)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011405144550415)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0440155104041515)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_A5Q),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h005500550f0f0f87)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f4b0f0f3333ffff)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_A5Q),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c555c5c53555353)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_B5Q),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_CQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffde00120012ffde)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h030500050c050f05)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa00ff)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_CQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h008affba008affba)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff01dd10ff02ee2)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_B5Q),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f4b33003300)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9900009999000099)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_C5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ff3ffffcffcffff)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_DQ),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_B5Q),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_DO6),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3f3c0c0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffe000e0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f01d2ed1e2)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_C5Q),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_CQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_DQ),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefaeefaeefaaa)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0cc00)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_BO5),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_DQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ee00ee00ee00)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa00ff300030)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaffaa00aaf0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.Q(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0099000f0099000f)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_C5Q),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f990f9999)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_C5Q),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55550055)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I2(1'b1),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccaac0aac0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a6a6a6a6)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_DLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f2f0f000020000)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_CQ),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haacfaa0faac0aa00)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa00faffc800c8)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_ALUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_C5Q),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefefffffefe)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_DLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_DQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0f00ff00f0ff0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50fa50ee44)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000cc55cc55)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_ALUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hecec2020ecec2020)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc50cc05cc50)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0a0f0a0f0a0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fa50ee44fa50)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550055ff000000)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_A5Q),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa00c0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_CLUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcac0c00055ffff)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33300000)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_DO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa03300330)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0eeeeee00)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00fc0c)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_CQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccfacc00ccfa)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc30ffffec20)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_DQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_B5Q),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_DO6),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc00aaaafc00)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa0000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbe00be0c0c0c0c)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.R(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f5a3333)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_DQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacaca0cccccc00)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888fff00000)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_DQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0e4a0ff00cc00)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff3c003c)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa0000)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafb0051aafb0051)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeeea40404440)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffe0ffff00e0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222f3c0f3c0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_A5Q),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54aa00fcfc0000)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0a0f0a0f0a0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_CO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_DO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f0fc0003000c)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f505f000fa0a)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba10ba10ba10ba10)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3a0a0fa0afa0a)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_DQ),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_CO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_DO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05500550)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05500550)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffdfffdf)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_D5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd8d8ffffd888)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e0e0e0f0f0f00)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aafcaa00)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_CLUT (
.I0(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0f0aaaa)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafcfc)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_DQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_DO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaffffa0a0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_DLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005050ff005050)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeaaaafcf0fcf0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_DO6),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0eeeeeeaa)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_DO6),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5a0ee44ee44)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d888d88888d888d)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000088a888a8)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00af00af8caf8caf)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_ALUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1f5b1b1a0e4a0a0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_CQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000cfafa0a0a)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffef00ff00ef)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_A5Q),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa99aa55aa55)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I5(CLBLM_R_X11Y123_SLICE_X15Y123_CO6),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaaccf0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000cfafa0a0a)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff300030ffaa00aa)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5544aaaa5544aaa8)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11bb11aa00aa00)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0fdf805000d08)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30330000f0fff0ff)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f1f0fff0f1f0fff)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e0fffffffff)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00004010bfef)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055ffff30003000)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.R(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.R(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000af00f000f100)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7500880077008800)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fe22222323)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfcf0a0f0a0f)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303030201030102)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_CLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_D5Q),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000040)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff33ff30)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_ALUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555fcfc0c0c)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffccffffffcc)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc33333131)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_BO6),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I2(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_DO6),
.I5(CLBLM_L_X12Y115_SLICE_X17Y115_BQ),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafa0a0afa0a0a)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_BQ),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00fe00ff)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I2(CLBLM_L_X12Y115_SLICE_X17Y115_DO6),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_BO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X17Y115_AO6),
.Q(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X17Y115_BO6),
.Q(CLBLM_L_X12Y115_SLICE_X17Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X17Y115_CO6),
.Q(CLBLM_L_X12Y115_SLICE_X17Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeeffffffee)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_DLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d580d580)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_L_X12Y115_SLICE_X17Y115_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeaafaa45400500)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y115_SLICE_X17Y115_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb8bb8888b8b8888)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y115_SLICE_X17Y115_CQ),
.I5(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X16Y116_AO6),
.Q(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X16Y116_BO6),
.Q(CLBLM_L_X12Y116_SLICE_X16Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.Q(CLBLM_L_X12Y116_SLICE_X16Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccccffccff)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.I4(1'b1),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_DO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d580d580)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_CO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055445544)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_BQ),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefafdf5cc00cc00)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_AO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_AO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_BO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_DO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_CO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8f008fff800080)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I5(CLBLM_L_X12Y116_SLICE_X16Y116_CQ),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_BO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20ff33ec20cc00)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_AO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_AO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_CO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaaffffccc0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_C5Q),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00fc0000)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeccdc33320010)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I5(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X16Y118_AO6),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X16Y118_BO6),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555f0f00000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffa50ea40)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_CO6),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X16Y119_AO6),
.Q(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X16Y119_BO6),
.Q(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X16Y119_CO6),
.Q(CLBLM_L_X12Y119_SLICE_X16Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y119_SLICE_X16Y119_DO6),
.Q(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888d8d8d8d8)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_DO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0054540000)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_CO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0dfd0dfc0cfc0c)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_BLUT (
.I0(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_BO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffecccfcccec)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_AO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_DO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_CO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_BO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fff00000eeee)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_DQ),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_CQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_CQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_CO5),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_DO5),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_AO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_BO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_CO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_DO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4170417013441344)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_DLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_C5Q),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_D5Q),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a4c00cc05000aaa)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_CLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_C5Q),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_CQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_DQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf707f000f606f000)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_BLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000dcdedcde)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_CO5),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X17Y120_AO6),
.Q(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.Q(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_DLUT (
.I0(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I1(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I2(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_CO6),
.I4(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200aa0000540000)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_CLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I5(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff4f004fff400040)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_BLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888bb88b8b8bb88)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.R(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f992f2200000000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_DLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h001fffff11111111)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300222233002222)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_BLUT (
.I0(CLBLM_R_X13Y121_SLICE_X19Y121_DO6),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.I4(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cf55555554)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_AO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_BO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4b5affff5a5a)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_DLUT (
.I0(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa0515faea)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_CLUT (
.I0(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I3(CLBLM_R_X13Y121_SLICE_X19Y121_DO6),
.I4(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0f5f005000500)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_BLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y121_SLICE_X17Y121_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c5c5c0c5c0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.I4(1'b1),
.I5(CLBLM_L_X12Y121_SLICE_X17Y121_CO6),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f5f5f5f5)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_DLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h02020202005f005f)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_CLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2333ffff0c0c0000)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_BLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcccdc11100010)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X17Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.Q(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000313300003122)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_DLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_CO5),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000055000000)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_CLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I1(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000fd0df808)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I1(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffffa200a2)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_ALUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_BO6),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I5(CLBLM_L_X12Y122_SLICE_X17Y122_CO6),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_BO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_CO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0aca00000aca)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_CLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1c0d1d1c0d1c0c0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22332233a2f3a2f3)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_DQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y123_SLICE_X15Y123_DO6),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_AO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_BO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000efff0000fdff)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_DLUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I4(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4f50f0ff0f0a0a0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_CLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505fd0df000f808)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I4(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333ff002121)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_DO6),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.R(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0000000aaaa0000)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_ALUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33335fff00005fff)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h23232323afafafaf)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa800080008000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f10101f4f40404)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_BQ),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeaeaccccc0c0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000eccca000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc00fff000f0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_A5Q),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y113_SLICE_X7Y113_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe0ffe0e0e0e0e0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_CQ),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0acc00cc0acc00)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h400040000fff0fff)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffef5545aaea0040)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I4(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcddc0110dcdc1010)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_DO6),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeccfefe32003232)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_DQ),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcdcdcd01010101)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_CQ),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff00fcfc0000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_BQ),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf3ffc000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaf69966996)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffc0cf505f404)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acacacaca)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffac80000fac8)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_BQ),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.Q(CLBLM_R_X3Y118_SLICE_X2Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8aaa8aaa8a8a8a8a)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h113355ffc33c3cc3)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f088882288)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_BQ),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20ce02ec20ce02)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_CQ),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabbabffffffff)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_A5Q),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_A5Q),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb0bf4f40b)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f0cccc)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aaf0aaf0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.Q(CLBLM_R_X3Y119_SLICE_X2Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.Q(CLBLM_R_X3Y119_SLICE_X2Y119_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.Q(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.Q(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0000070f0800)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_BQ),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_A5Q),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_B5Q),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f88888fffff00ff)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_B5Q),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_A5Q),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ffaaaaaa)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaacccc)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_DQ),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3bff33ff3fff33)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aa30aaffaa00)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_CQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0c0c0c0c)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_CQ),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf5f5a0a0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.Q(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f0f0f55550000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I3(1'b1),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff30ffba3030baba)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcccdccc5000dccc)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0ccf0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_DQ),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.Q(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.Q(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.Q(CLBLM_R_X3Y120_SLICE_X3Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000033000a0a3b0a)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I3(LIOB33_X0Y65_IOB_X0Y66_I),
.I4(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0c5c00000c5c)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20cc00cc00cc00)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_BQ),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_A5Q),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdec3120ffcc3300)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_BQ),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111000055115500)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22002200aaaa2200)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I2(1'b1),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_B5Q),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3b0a3b0a)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_DQ),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I3(LIOB33_X0Y63_IOB_X0Y63_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffa)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_BO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.Q(CLBLM_R_X3Y121_SLICE_X3Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.Q(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7755330077553300)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.I2(1'b1),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50dcffff50dc50dc)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I3(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(CLBLL_L_X2Y124_SLICE_X1Y124_CO6),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_CO6),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_DO6),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fa50ee44fa50)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_A5Q),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040455045504)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I1(LIOB33_X0Y71_IOB_X0Y71_I),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_DQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff30baffff30ba)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.I2(LIOB33_X0Y67_IOB_X0Y67_I),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00000ace0a0a)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y67_I),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffffffdfff)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff2f2fffff2222)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.I3(1'b1),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff30baffff30ba)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_CQ),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafaaaaefefeeee)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_CO6),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeffffffffffefff)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff50dc50dc)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_CQ),
.I2(LIOB33_X0Y53_IOB_X0Y54_I),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_BO6),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdfcfdfc)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_AO6),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AO6),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccdddc00001110)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_A5Q),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbfffffffa)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_CO6),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_BO6),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_BO6),
.I4(CLBLM_R_X5Y123_SLICE_X6Y123_BO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_CQ),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceefcfe00aaf0fa)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_A5Q),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I2(LIOB33_X0Y65_IOB_X0Y65_I),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefffe)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_DO6),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_DO6),
.I3(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.I4(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_DO6),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f4fff4f4444ff44)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_AO6),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_DQ),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000044440f004f44)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_DQ),
.I4(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000f000000080)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_DLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_AO6),
.I5(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcfdfcfcfc)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_CLUT (
.I0(CLBLM_R_X3Y125_SLICE_X2Y125_AO6),
.I1(CLBLL_L_X2Y124_SLICE_X1Y124_BO6),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_DO6),
.I5(CLBLL_L_X2Y124_SLICE_X0Y124_CO6),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_BLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_BO6),
.I1(CLBLL_L_X2Y124_SLICE_X1Y124_CO6),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_CO6),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefefffffffe)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_ALUT (
.I0(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_DO6),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_CO6),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I4(CLBLL_L_X2Y124_SLICE_X0Y124_BO6),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff22fff2)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_DLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_DQ),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_CO6),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I5(CLBLM_R_X5Y122_SLICE_X7Y122_DO6),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff111f11ff000f00)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_CLUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_CQ),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333233100000050)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7ffffffdf)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdfffffffff)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0c00aa0cae)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_DQ),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I2(CLBLM_R_X3Y126_SLICE_X2Y126_BO6),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_AO5),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_DO6),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_AO6),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_BLUT (
.I0(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_CO6),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_BO6),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_AO6),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0000000afafffff)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff700000400)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffffffffffff)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000eeecaaa0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfff5fff00008000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h52555a5588000000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000faf80a08)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff210000002100)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_DQ),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05000500aaee0044)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaabe00fc003c)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cf000f000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f40004fbfbfbfb)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffffffffffff)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_CQ),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4f5e4f5e4a0a0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808f808fc0cfc0c)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001212ff003030)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_BO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_CO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_DO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888ddd88888)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_DQ),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_CQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ee44ee44)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_C5Q),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f30003f0fc000c)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88d888ff00f000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf000aaaa3c00)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_DQ),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01144f0f01144)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808ff0ff808f000)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aaccaac0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_C5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333303333)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffefee)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccffcc00)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00c8000000c8)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000005000cc00cc)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54aa00fe54fe54)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fafaff00c8c8)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccccccffc0c0c0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1c081f0f0c0c0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1a081f0f0a0a0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f0f003030000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f60006f0f60006)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_BO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c033773377)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc00fc00ff00aa00)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_A5Q),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cccc5a5a)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f505fa0a)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_DQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffdfffffffffff)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22ed21ed21)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ccccefcf)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000faf8f0f8)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffaa)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4a0e4f5e4a0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaffeaee50554044)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00cc00c0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X7Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff5)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_B5Q),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_D5Q),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff02)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff505050505050)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_CO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffffff)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fff0f03300)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_DQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_C5Q),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0cfc0c0cfc0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888d888d888)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccffccffcc)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_D5Q),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_B5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc55f0cccc00f0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_DQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000b8aab8aa)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_C5Q),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf000f0cc)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ff0000f00000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff000404)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000000000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000010000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_CQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_A5Q),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f00aaaacccc)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333cece0202)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_CO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001000000010)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_DLUT (
.I0(CLBLM_R_X29Y141_SLICE_X42Y141_AO6),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heccccccc20000000)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_CLUT (
.I0(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0cccc)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00fcfc)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7733550077335500)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.I2(1'b1),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1055101010551010)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_CLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0caaffaacc)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff00fdfd)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00afaaafaa)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_DLUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000005400000010)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_CLUT (
.I0(CLBLM_R_X29Y141_SLICE_X42Y141_AO6),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0afacacacac)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555000005550)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_ALUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_CO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111000051515050)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_DLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaefeae54045404)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_D5Q),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f0ffcc)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e2e2ff00aaaa)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_ALUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CQ),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505040401010000)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_DLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.I3(1'b1),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000000ca)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLM_R_X29Y141_SLICE_X42Y141_AO6),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002200000030)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_BLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_DQ),
.I1(CLBLM_R_X29Y141_SLICE_X42Y141_AO6),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff77fffffffffb)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_BO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_CO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaaeeffffaaee)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_CQ),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00ee44ee44)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00cccc)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaf00000aaf0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_ALUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_AO5),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_CO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1013101000030000)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_CLUT (
.I0(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_DQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00440f4f00440044)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_BLUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I2(CLBLL_L_X2Y123_SLICE_X1Y123_DO6),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.I4(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfff0ff00)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ffaa5500)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_DQ),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeaaaea00400040)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404f404f404)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff004800000048)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550055ff500050)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00066f0f00000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_C5Q),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f8f8f822888888)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff282828ffa0a0a0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf088880000)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_CLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(RIOB33_X105Y127_IOB_X1Y127_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf222f888f222f888)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f8f4f844884488)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_ALUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_CO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaac000c000)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0b1a011001100)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000202ff002020)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y126_SLICE_X5Y126_AO6),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0a0a0e4a0a0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d88d888888888)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.Q(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.Q(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05544f0f00000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaa3030)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_DQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020200000202)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0e4a0e4a0e4)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_B5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0f04444)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff00a8a8)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000505)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafffee00000000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DQ),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0efe0ef000f000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_A5Q),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccff00)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff0000af0000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3310333333103333)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff000ff0fc000c)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0002020000fafa)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50fe54ba10)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_DQ),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_DO6),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4a0000000ff)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_B5Q),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003232ff000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffefffffff)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.I2(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0ccf0cc)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_A5Q),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf80d08f5f00500)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fe10fe10)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaf0505aeae0404)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0dd88f0f05500)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fff0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_DQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888dddd8888)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff55aa00aa00)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0cac0c5c0ca)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeaaba55540010)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_AQ),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffc)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_B5Q),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_C5Q),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54aa00aa00)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_CQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0010101010)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_D5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0afc0cf000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc000f00f0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_A5Q),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a0a3a0aca0ac)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f101f404f404)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeec0cceeeaccc0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1212212184844848)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a2a080808080)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff10efffffdddd)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ff5000500050)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000fffe)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_DLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_DO6),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.I4(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0506050505050505)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_CQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f6ac06ac0953f95)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.I4(CLBLM_L_X12Y119_SLICE_X16Y119_DQ),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0af606fa0afa0a)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_CLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.I4(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cfcfcfcac0c0c0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_BLUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05050505f5f5f5f5)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd01cc00aaaa0000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_DO6),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003030aaaaff0f)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0aca0accfcfc0c0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc55f5cccc00f0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_CO6),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff00fc)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_A5Q),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcccece30303030)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000f0f0c0c)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd8ddd88888)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33cc3c33cc33c)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_A5Q),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fc00fc00ff00aa)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_A5Q),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaaaaaf8f88888)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f0f6f006000600)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_DQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3133313331331133)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefffeff0f000f00)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafacaca0a0acac)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_DQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_A5Q),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfd0d0df1fd010d)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff7)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb111100cf00cf)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafaee50505044)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00fa05050505)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffbfff)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00e0e0e0e0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_A5Q),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe0e0ef4f40404)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fcaaaa00fc)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fd00fd00fd00)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5e4a0a0f5e4)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f50505f4f40404)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbaafaaa51005000)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaabbaa11001100)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0b1b1b1b1a0a0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff30f03fcf00c00)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00f000f000f0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_CO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_DO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ff55aa00)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044d8d8d8d8)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555f0f04444)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5550cccc5550)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_ALUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_DO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8bb88b8b8bb88)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_DLUT (
.I0(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_DQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5e4a0a0f5e4)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_CQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_CQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_D5Q),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff0c0ffcf00c00)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaf0aaf0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_CQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff15ff3f80800000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_CLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_DO6),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6fc66ccf0f00000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_A5Q),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hde5afcf0cc00cc00)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_ALUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_CO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_DO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd888d888d8)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_CQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_DQ),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ee44ef45)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_A5Q),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff6fff60f060f06)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_BLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_DO6),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdc505033003300)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f1f5f3fff3fff)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3cbe3caa00aa00)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000fcfc3030)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff000ff0f00000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000aa000000aa)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habaeaeae01040404)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfc0cfc0c0c0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f80808f4f80408)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f60006f0f00000)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff00f0f0f00)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_BQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_B5Q),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa50fa50)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_ALUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555655ff33ff33)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_DQ),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfddd3111eccc2000)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_CO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000fa500003333)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_DLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaeeaa55004400)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfcfa0c0a)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_BLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff10effdfdfdfd)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_DQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X15Y114_AO6),
.Q(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.Q(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcf0f00f0c0000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(CLBLM_L_X12Y116_SLICE_X16Y116_CQ),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc50cc00cc00)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X12Y115_SLICE_X17Y115_BQ),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d7d7dbebebebe)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699669966996)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011223302132031)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_B5Q),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002200f0f0e1f0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_CO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cffff3c3cffff3c)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5fafffff5fa)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_DO6),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_CQ),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I2(CLBLM_L_X12Y115_SLICE_X17Y115_CQ),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I5(CLBLM_L_X12Y116_SLICE_X16Y116_CQ),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5fdf5f5f5f7f)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_CO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_CO6),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_BO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2112122121121221)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0fff088f0cc)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0aa00aaff)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_DQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550055ff500050)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I5(CLBLM_L_X12Y116_SLICE_X16Y116_BQ),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6f6f6ff6f6f6f6)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_DLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff6ff6ffff6ff6)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f0f0f3fff0f0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffabff03aaaa0000)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2323232301010101)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000cfcf)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_DQ),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fafa0a0a)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_CQ),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_D5Q),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fcfc0000)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_BO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_CO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb8ffb8ffb8ff88)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_DQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccaa00aa)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c0c0ff00aaaa)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc50050000)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_BO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002200000002)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_DLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cccc000a000a)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff6fff60f060f06)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_DO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_CQ),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000445500)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_ALUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_DO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22ec20ec20)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_DQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaab0001aaae0004)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c0c0aaaa)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff51ff5100510051)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_BQ),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_BO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_CO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaafaeafaea)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_DO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaa05000500)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00e0e0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_BQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00f000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_DQ),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heccccccca0000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_DLUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020202002222222)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_CLUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0010104040)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_BLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8a8a8ffa0a0a0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_ALUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_DLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_DO6),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcfc00)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0a0acccc0a0a)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_DQ),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aaffaaf0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_CO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_DO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaaaa55540000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff55aa00ab01)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0aca00000aca)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_DQ),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccedcccc00210000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_CQ),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080008000000)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f202f202f000)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_A5Q),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffac00aa00ac)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_BLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00fc30)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_ALUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_CO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffccc4c4ffc4)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_DLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_CO6),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeaa44554400)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I5(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404ff0ff404f000)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_BLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ee4405050000)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_CQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_BO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_CO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500ccccf5a0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_DLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaa00fc)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_CLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I3(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0205010ff33ff33)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_BLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefff0000efff)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_DQ),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0acccc0000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_DLUT (
.I0(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h72325f1fddddf0f0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000660033)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_CO6),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7077303370773033)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_ALUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_BO6),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.R(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0000000c0c0c0c)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_DLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_AO6),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3031323333333333)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_CLUT (
.I0(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_AO6),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3000cfff2000df)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_BLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_AO6),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.I4(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200220022)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_ALUT (
.I0(CLBLM_R_X11Y122_SLICE_X15Y122_DO6),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5aaa59aa55aa55)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_DLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.I4(CLBLM_R_X11Y122_SLICE_X15Y122_DO6),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5070000000000a08)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff737f)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_BLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_DO6),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010101000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h99999999aa99a999)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I4(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3313333333333323)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_CLUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h40cc50ff40cc50ff)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_BLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_DO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf33f333351151111)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_BO6),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X15Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h404040c000000000)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_B5Q),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h99ff00ff090f000f)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_BLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_CO6),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f4f4ff00f4f4)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf03cf03cf00ff00f)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22a233f322a233f3)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_ALUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_DQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0fcf0fc)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b888b88aaaaffff)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_ALUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y115_SLICE_X18Y115_AO6),
.Q(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y115_SLICE_X18Y115_BO6),
.Q(CLBLM_R_X13Y115_SLICE_X18Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_DO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_CO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccfcccfc)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_B5Q),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_BQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_BO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0cca0cc00ccff)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_BQ),
.I2(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_BO6),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_AO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_DO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_CO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_BO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_AO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y120_SLICE_X18Y120_AO6),
.Q(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y120_SLICE_X18Y120_BO6),
.Q(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005040000)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_DLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I3(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a2a000000000000)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_CLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I5(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_CO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5f5f5a0)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_AQ),
.I3(CLBLM_R_X13Y121_SLICE_X19Y121_AO6),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_BO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcdddc11101110)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.I3(CLBLM_R_X13Y121_SLICE_X19Y121_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y119_SLICE_X16Y119_CQ),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_AO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_DO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_CO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000030000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I4(CLBLM_R_X13Y120_SLICE_X18Y120_DO6),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_BO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ffffffffffffff)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_ALUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_CO6),
.I1(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I4(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_AO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y121_SLICE_X18Y121_AO6),
.Q(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y121_SLICE_X18Y121_BO6),
.Q(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333fffffff7)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_DLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_DO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000dfdfcfff)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_CLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_CO6),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_BQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_DO6),
.I4(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_CO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0bff0e000b000e)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_BLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.I1(CLBLM_R_X13Y121_SLICE_X19Y121_BO6),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CQ),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_BO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccfacc00ccaf)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_ALUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_CO6),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_AO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_DLUT (
.I0(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I1(CLBLM_R_X13Y120_SLICE_X18Y120_DO6),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I4(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_BQ),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_DO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0ff5f00e0ff1f0)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_CLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I1(CLBLM_R_X13Y120_SLICE_X19Y120_AO6),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_BQ),
.I4(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I5(CLBLM_R_X13Y120_SLICE_X19Y120_BO6),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_CO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccdccccccefcccc)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_BLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I2(CLBLM_R_X13Y122_SLICE_X19Y122_AO6),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I5(CLBLM_R_X13Y122_SLICE_X19Y122_BO6),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_BO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c2d3c0f3c3c3c3c)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_ALUT (
.I0(CLBLM_R_X13Y122_SLICE_X19Y122_BO6),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I2(CLBLM_R_X13Y120_SLICE_X18Y120_BQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I4(CLBLM_R_X13Y122_SLICE_X19Y122_AO6),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_AO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X18Y122_AO6),
.Q(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y122_SLICE_X18Y122_BO6),
.Q(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5fafaf5f5f5fa)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_DLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I4(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_DO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100001000)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_CLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_CO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202f202f202f202)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_BLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_DO6),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_BO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfc3130fdfc3130)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_AO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_DO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_CO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffffff)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_BLUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I4(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_BO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.I2(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I3(CLBLM_L_X12Y121_SLICE_X17Y121_BQ),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_AO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33c933cc33c633cc)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_CLUT (
.I0(CLBLM_R_X13Y122_SLICE_X18Y122_BQ),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_CQ),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30300005cf45aa50)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_BLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I3(CLBLM_L_X12Y120_SLICE_X16Y120_BQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff0ffa0a)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_ALUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_CO6),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y141_SLICE_X42Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y141_SLICE_X42Y141_DO5),
.O6(CLBLM_R_X29Y141_SLICE_X42Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y141_SLICE_X42Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y141_SLICE_X42Y141_CO5),
.O6(CLBLM_R_X29Y141_SLICE_X42Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y141_SLICE_X42Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y141_SLICE_X42Y141_BO5),
.O6(CLBLM_R_X29Y141_SLICE_X42Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbfbfbfffffafa)
  ) CLBLM_R_X29Y141_SLICE_X42Y141_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(1'b1),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLM_R_X29Y141_SLICE_X42Y141_AO5),
.O6(CLBLM_R_X29Y141_SLICE_X42Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y141_SLICE_X43Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y141_SLICE_X43Y141_DO5),
.O6(CLBLM_R_X29Y141_SLICE_X43Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y141_SLICE_X43Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y141_SLICE_X43Y141_CO5),
.O6(CLBLM_R_X29Y141_SLICE_X43Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y141_SLICE_X43Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y141_SLICE_X43Y141_BO5),
.O6(CLBLM_R_X29Y141_SLICE_X43Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y141_SLICE_X43Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y141_SLICE_X43Y141_AO5),
.O6(CLBLM_R_X29Y141_SLICE_X43Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_DO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_CO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_BO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202020202020202)
  ) CLBLM_R_X37Y120_SLICE_X56Y120_ALUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X56Y120_AO5),
.O6(CLBLM_R_X37Y120_SLICE_X56Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_DO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_CO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_BO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y120_SLICE_X57Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y120_SLICE_X57Y120_AO5),
.O6(CLBLM_R_X37Y120_SLICE_X57Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_ALUT (
.I0(RIOB33_X105Y139_IOB_X1Y139_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffff0f0ffff)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffccffccff)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33f3f3f3f3)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ffccffccff)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I2(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_BO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_BO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_CO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X8Y124_SLICE_X10Y124_DQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X4Y118_SLICE_X4Y118_CQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y124_SLICE_X10Y124_D5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X5Y115_SLICE_X7Y115_B5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X3Y117_SLICE_X3Y117_B5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X12Y123_D5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X3Y115_A5Q),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X5Y125_SLICE_X6Y125_CQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y138_SLICE_X163Y138_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X37Y120_SLICE_X56Y120_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_L_X12Y119_SLICE_X17Y119_AO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X10Y121_SLICE_X13Y121_DO6),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_L_X12Y119_SLICE_X17Y119_AO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X10Y121_SLICE_X13Y121_DO6),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X12Y119_SLICE_X16Y119_BQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_R_X11Y124_SLICE_X15Y124_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y115_SLICE_X18Y115_BQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X29Y141_SLICE_X42Y141_AO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X29Y141_SLICE_X42Y141_AO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_AMUX = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_BMUX = CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_AMUX = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_BMUX = CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_CMUX = CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_BMUX = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AMUX = CLBLL_L_X2Y119_SLICE_X1Y119_A5Q;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_BMUX = CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_BMUX = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_AMUX = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_AMUX = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_BMUX = CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_CMUX = CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_AMUX = CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B = CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_AMUX = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B = CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D = CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D = CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_AMUX = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_AMUX = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_BMUX = CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_DMUX = CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_DMUX = CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_CMUX = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_DMUX = CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CMUX = CLBLL_L_X4Y118_SLICE_X4Y118_C5Q;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_AMUX = CLBLL_L_X4Y119_SLICE_X4Y119_A5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CMUX = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_CMUX = CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_DMUX = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_AMUX = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_AMUX = CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A = CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B = CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A = CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_BMUX = CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A = CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_AMUX = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_CMUX = CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_AMUX = CLBLM_L_X8Y113_SLICE_X10Y113_A5Q;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_BMUX = CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_BMUX = CLBLM_L_X8Y113_SLICE_X11Y113_B5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_AMUX = CLBLM_L_X8Y114_SLICE_X11Y114_A5Q;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_BMUX = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_AMUX = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_BMUX = CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_DMUX = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_BMUX = CLBLM_L_X8Y116_SLICE_X11Y116_B5Q;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A = CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B = CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CMUX = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_CMUX = CLBLM_L_X8Y117_SLICE_X11Y117_C5Q;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_BMUX = CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_DMUX = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_AMUX = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CMUX = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_DMUX = CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CMUX = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_BMUX = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_DMUX = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_AMUX = CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_BMUX = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A = CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_AMUX = CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CMUX = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_DMUX = CLBLM_L_X8Y123_SLICE_X10Y123_D5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CMUX = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A = CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B = CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CMUX = CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_DMUX = CLBLM_L_X8Y124_SLICE_X10Y124_D5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A = CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_AMUX = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CMUX = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A = CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CMUX = CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_DMUX = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A = CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_DMUX = CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A = CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_AMUX = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_BMUX = CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_AMUX = CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_BMUX = CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_CMUX = CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_DMUX = CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_AMUX = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_BMUX = CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_DMUX = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_AMUX = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_CMUX = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B = CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_BMUX = CLBLM_L_X10Y115_SLICE_X12Y115_B5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_CMUX = CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_AMUX = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_BMUX = CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_AMUX = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_BMUX = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_AMUX = CLBLM_L_X10Y118_SLICE_X12Y118_A5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_AMUX = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_AMUX = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_BMUX = CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CMUX = CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_AMUX = CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_BMUX = CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CMUX = CLBLM_L_X10Y120_SLICE_X12Y120_C5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_DMUX = CLBLM_L_X10Y120_SLICE_X12Y120_D5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_AMUX = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_DMUX = CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_AMUX = CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_BMUX = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_DMUX = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_DMUX = CLBLM_L_X10Y122_SLICE_X13Y122_D5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_DMUX = CLBLM_L_X10Y123_SLICE_X12Y123_D5Q;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_DMUX = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_AMUX = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_AMUX = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_BMUX = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A = CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_BMUX = CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B = CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A = CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A = CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B = CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A = CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B = CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D = CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A = CLBLM_L_X12Y116_SLICE_X17Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B = CLBLM_L_X12Y116_SLICE_X17Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C = CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D = CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A = CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B = CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A = CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C = CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D = CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A = CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B = CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C = CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A = CLBLM_L_X12Y119_SLICE_X16Y119_AO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B = CLBLM_L_X12Y119_SLICE_X16Y119_BO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C = CLBLM_L_X12Y119_SLICE_X16Y119_CO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D = CLBLM_L_X12Y119_SLICE_X16Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B = CLBLM_L_X12Y119_SLICE_X17Y119_BO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C = CLBLM_L_X12Y119_SLICE_X17Y119_CO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_AMUX = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B = CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C = CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D = CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_CMUX = CLBLM_L_X12Y120_SLICE_X16Y120_C5Q;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_DMUX = CLBLM_L_X12Y120_SLICE_X16Y120_D5Q;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A = CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_AMUX = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_BMUX = CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_CMUX = CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A = CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B = CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_DMUX = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A = CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_BMUX = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_CMUX = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_DMUX = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A = CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_CMUX = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B = CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A = CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B = CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_CMUX = CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_AMUX = CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A = CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B = CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C = CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AMUX = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CMUX = CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_CMUX = CLBLM_R_X3Y116_SLICE_X2Y116_C5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_DMUX = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_CMUX = CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_BMUX = CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_DMUX = CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_CMUX = CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_CMUX = CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_AMUX = CLBLM_R_X3Y119_SLICE_X2Y119_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_BMUX = CLBLM_R_X3Y119_SLICE_X2Y119_B5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_CMUX = CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_DMUX = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_AMUX = CLBLM_R_X3Y121_SLICE_X3Y121_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_AMUX = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_AMUX = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_AMUX = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_DMUX = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_AMUX = CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_BMUX = CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_CMUX = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_AMUX = CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_AMUX = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_CMUX = CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_DMUX = CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_AMUX = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_BMUX = CLBLM_R_X5Y113_SLICE_X7Y113_B5Q;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_DMUX = CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_AMUX = CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_BMUX = CLBLM_R_X5Y115_SLICE_X7Y115_B5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_DMUX = CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CMUX = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CMUX = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_DMUX = CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CMUX = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CMUX = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CMUX = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_BMUX = CLBLM_R_X5Y120_SLICE_X7Y120_B5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A = CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B = CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C = CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_AMUX = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A = CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B = CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C = CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A = CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_AMUX = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A = CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A = CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_CMUX = CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AMUX = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_BMUX = CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CMUX = CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CMUX = CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_AMUX = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_BMUX = CLBLM_R_X7Y114_SLICE_X8Y114_B5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_BMUX = CLBLM_R_X7Y114_SLICE_X9Y114_B5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_CMUX = CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_CMUX = CLBLM_R_X7Y115_SLICE_X8Y115_C5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_AMUX = CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_AMUX = CLBLM_R_X7Y116_SLICE_X9Y116_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_BMUX = CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_AMUX = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_CMUX = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_DMUX = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_BMUX = CLBLM_R_X7Y119_SLICE_X8Y119_B5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CMUX = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_DMUX = CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_AMUX = CLBLM_R_X7Y119_SLICE_X9Y119_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CMUX = CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CMUX = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CMUX = CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_AMUX = CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CMUX = CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_AMUX = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CMUX = CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_DMUX = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_DMUX = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A = CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B = CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CMUX = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_DMUX = CLBLM_R_X7Y123_SLICE_X8Y123_D5Q;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A = CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B = CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CMUX = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A = CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B = CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_AMUX = CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_DMUX = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_BMUX = CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_AMUX = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_AMUX = CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_AMUX = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_CMUX = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_BMUX = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A = CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A = CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B = CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_CMUX = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_DMUX = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A = CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_CMUX = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_DMUX = CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A = CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_AMUX = CLBLM_R_X11Y121_SLICE_X14Y121_A5Q;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_AMUX = CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_DMUX = CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_AMUX = CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A = CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A = CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A = CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A = CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B = CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_AMUX = CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A = CLBLM_R_X13Y115_SLICE_X18Y115_AO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B = CLBLM_R_X13Y115_SLICE_X18Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C = CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D = CLBLM_R_X13Y115_SLICE_X18Y115_DO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A = CLBLM_R_X13Y115_SLICE_X19Y115_AO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B = CLBLM_R_X13Y115_SLICE_X19Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C = CLBLM_R_X13Y115_SLICE_X19Y115_CO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D = CLBLM_R_X13Y115_SLICE_X19Y115_DO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A = CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B = CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A = CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B = CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C = CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D = CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_AMUX = CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A = CLBLM_R_X13Y121_SLICE_X18Y121_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B = CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C = CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_DMUX = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A = CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B = CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C = CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D = CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A = CLBLM_R_X13Y122_SLICE_X18Y122_AO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B = CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_CMUX = CLBLM_R_X13Y122_SLICE_X18Y122_CO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A = CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B = CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C = CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A = CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B = CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_BMUX = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_CMUX = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A = CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B = CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C = CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D = CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_A = CLBLM_R_X29Y141_SLICE_X42Y141_AO6;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_B = CLBLM_R_X29Y141_SLICE_X42Y141_BO6;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_C = CLBLM_R_X29Y141_SLICE_X42Y141_CO6;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_D = CLBLM_R_X29Y141_SLICE_X42Y141_DO6;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_AMUX = CLBLM_R_X29Y141_SLICE_X42Y141_AO5;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_A = CLBLM_R_X29Y141_SLICE_X43Y141_AO6;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_B = CLBLM_R_X29Y141_SLICE_X43Y141_BO6;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_C = CLBLM_R_X29Y141_SLICE_X43Y141_CO6;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_D = CLBLM_R_X29Y141_SLICE_X43Y141_DO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B = CLBLM_R_X37Y120_SLICE_X56Y120_BO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C = CLBLM_R_X37Y120_SLICE_X56Y120_CO6;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D = CLBLM_R_X37Y120_SLICE_X56Y120_DO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A = CLBLM_R_X37Y120_SLICE_X57Y120_AO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B = CLBLM_R_X37Y120_SLICE_X57Y120_BO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C = CLBLM_R_X37Y120_SLICE_X57Y120_CO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D = CLBLM_R_X37Y120_SLICE_X57Y120_DO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A = CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B = CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C = CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D = CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B = CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C = CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D = CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_AMUX = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A = CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B = CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C = CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D = CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B = CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C = CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D = CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_AMUX = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y124_SLICE_X10Y124_D5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X5Y115_SLICE_X7Y115_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X10Y123_SLICE_X12Y123_D5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X29Y141_SLICE_X42Y141_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X29Y141_SLICE_X42Y141_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = CLBLM_R_X3Y119_SLICE_X3Y119_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = CLBLM_R_X3Y119_SLICE_X3Y119_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = CLBLM_R_X3Y117_SLICE_X2Y117_DQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_AX = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = CLBLM_R_X5Y120_SLICE_X7Y120_B5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = CLBLM_R_X3Y118_SLICE_X2Y118_BQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = CLBLM_R_X3Y119_SLICE_X2Y119_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = CLBLM_R_X3Y119_SLICE_X2Y119_B5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B6 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D3 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_B5Q;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = CLBLM_R_X3Y118_SLICE_X2Y118_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = CLBLM_R_X3Y119_SLICE_X2Y119_A5Q;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = CLBLM_R_X3Y120_SLICE_X3Y120_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = CLBLL_L_X4Y118_SLICE_X5Y118_DQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A1 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A3 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A5 = CLBLM_L_X12Y115_SLICE_X17Y115_CQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A6 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B2 = CLBLM_L_X12Y115_SLICE_X17Y115_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B4 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C2 = CLBLM_L_X12Y115_SLICE_X17Y115_CQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C5 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D1 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D2 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D5 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D6 = 1'b1;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C6 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A2 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A3 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A4 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A5 = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A6 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B1 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B3 = CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B4 = CLBLM_L_X12Y115_SLICE_X17Y115_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B5 = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B6 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C1 = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C2 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C3 = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C5 = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C6 = CLBLM_L_X12Y115_SLICE_X17Y115_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D2 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D4 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = CLBLM_R_X3Y119_SLICE_X2Y119_A5Q;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_AX = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A6 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = CLBLM_R_X3Y117_SLICE_X2Y117_DQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = CLBLM_R_X3Y119_SLICE_X2Y119_B5Q;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A3 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A4 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A6 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B2 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B5 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B6 = CLBLM_L_X12Y116_SLICE_X16Y116_CQ;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C4 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_A6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D4 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A1 = CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A3 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A4 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A6 = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C2 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B1 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B2 = CLBLM_L_X12Y116_SLICE_X16Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B3 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B4 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C2 = CLBLM_L_X12Y116_SLICE_X16Y116_CQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C5 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_A6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D2 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D3 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D4 = CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D5 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D6 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_C6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D1 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D2 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D3 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D5 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = CLBLM_R_X3Y117_SLICE_X3Y117_CQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = CLBLM_R_X5Y115_SLICE_X6Y115_DQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A4 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B4 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C4 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D4 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A3 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A5 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A6 = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = CLBLM_R_X5Y115_SLICE_X7Y115_B5Q;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B1 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B2 = CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B3 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C1 = CLBLM_R_X3Y116_SLICE_X2Y116_C5Q;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C2 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C5 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D4 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_AX = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_B5Q;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = CLBLM_R_X5Y125_SLICE_X6Y125_DQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = CLBLM_R_X5Y125_SLICE_X6Y125_DQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = CLBLM_R_X3Y120_SLICE_X3Y120_CQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = CLBLM_R_X3Y121_SLICE_X3Y121_A5Q;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = CLBLM_R_X3Y120_SLICE_X3Y120_CQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A3 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A4 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A6 = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B3 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_B5Q;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A4 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B5 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C1 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C2 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C4 = CLBLL_L_X4Y116_SLICE_X4Y116_CQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C6 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D2 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D3 = CLBLM_R_X7Y124_SLICE_X9Y124_DQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D4 = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D5 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D6 = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A1 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A2 = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A3 = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A4 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A5 = CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A6 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B1 = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B2 = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B3 = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B4 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B5 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B6 = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C1 = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C2 = CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C3 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C4 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C5 = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C6 = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D1 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D2 = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D3 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D5 = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A1 = CLBLM_L_X10Y118_SLICE_X13Y118_DQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A2 = CLBLM_L_X12Y119_SLICE_X16Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A4 = CLBLM_L_X12Y117_SLICE_X16Y117_CQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A6 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B1 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B2 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B3 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B4 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B6 = 1'b1;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C1 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C2 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C3 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C4 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D1 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D2 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D3 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D4 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D6 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A2 = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A3 = CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A6 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B1 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B2 = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B4 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C2 = CLBLM_L_X12Y119_SLICE_X16Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C3 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D2 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D3 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D4 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A1 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D3 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B2 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = CLBLM_R_X3Y119_SLICE_X3Y119_CQ;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D6 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D6 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C5 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B1 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B2 = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B4 = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B5 = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B6 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C1 = CLBLM_R_X7Y124_SLICE_X9Y124_DQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C2 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C3 = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C4 = CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C5 = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C6 = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D3 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A1 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A3 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A4 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A5 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A6 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B1 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B2 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B3 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B6 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C1 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C2 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C3 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C4 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C5 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C6 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D1 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D2 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D3 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D4 = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D5 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D6 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A1 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A2 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A4 = CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A5 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B1 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B2 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B6 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B4 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C1 = CLBLM_L_X12Y120_SLICE_X16Y120_C5Q;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C3 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C5 = CLBLM_L_X12Y120_SLICE_X16Y120_D5Q;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D1 = CLBLM_L_X12Y120_SLICE_X16Y120_C5Q;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D2 = CLBLM_L_X12Y120_SLICE_X16Y120_D5Q;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D3 = CLBLM_L_X12Y120_SLICE_X16Y120_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B5 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D5 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C2 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C3 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C4 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C2 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D2 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X29Y141_SLICE_X42Y141_AO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C6 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X29Y141_SLICE_X42Y141_AO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A1 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A2 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A4 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A6 = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B1 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B4 = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B6 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C1 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C2 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C3 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C4 = CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C5 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C6 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D1 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D2 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D3 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D4 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D5 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D6 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A1 = CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A2 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A4 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A5 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_C6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_AX = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B1 = CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B2 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B4 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B5 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C4 = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C5 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D2 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D3 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D4 = CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D5 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D6 = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_SR = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A2 = CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A3 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A5 = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A6 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B1 = CLBLM_L_X8Y113_SLICE_X11Y113_B5Q;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B2 = CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B4 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A1 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A2 = CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A3 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A5 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A6 = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B2 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B4 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B5 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B6 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = CLBLM_L_X8Y113_SLICE_X10Y113_A5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C1 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C2 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C3 = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D1 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_A5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D6 = CLBLM_R_X13Y122_SLICE_X18Y122_CO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D4 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A5 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A6 = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B1 = CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B2 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B3 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B4 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B5 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C1 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C2 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C3 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A5 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B1 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B5 = CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C1 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C4 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C5 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D1 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A1 = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A3 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A4 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A6 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B2 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B5 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B6 = CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C1 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D5 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D6 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = CLBLM_L_X8Y113_SLICE_X11Y113_B5Q;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D4 = CLBLM_L_X12Y123_SLICE_X17Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A1 = CLBLM_R_X11Y117_SLICE_X15Y117_DQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A3 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A5 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A6 = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B3 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B4 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B5 = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = CLBLM_L_X12Y115_SLICE_X17Y115_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C1 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C2 = CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C3 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = CLBLM_R_X7Y114_SLICE_X9Y114_B5Q;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = CLBLM_R_X7Y116_SLICE_X9Y116_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C3 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C1 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C2 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C4 = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A4 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A5 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A6 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C5 = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A4 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C6 = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B4 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D3 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = CLBLM_R_X7Y116_SLICE_X9Y116_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = CLBLM_R_X5Y114_SLICE_X7Y114_DQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D5 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A3 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A4 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A1 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_C5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C4 = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C5 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_AX = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D2 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = CLBLM_R_X11Y118_SLICE_X15Y118_DQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = CLBLM_R_X7Y114_SLICE_X9Y114_B5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_SR = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = CLBLM_R_X7Y115_SLICE_X8Y115_C5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B4 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C4 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C5 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A2 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A4 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A1 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A3 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A6 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B1 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B2 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B3 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B5 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C1 = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C2 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C3 = CLBLM_R_X7Y115_SLICE_X8Y115_C5Q;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C5 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D3 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B5 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D1 = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D2 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D3 = CLBLM_R_X7Y115_SLICE_X8Y115_C5Q;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D4 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A1 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A2 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A5 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B5 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D1 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D2 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D4 = CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D5 = CLBLM_R_X11Y118_SLICE_X15Y118_DQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A4 = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B6 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C2 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C3 = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C4 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D5 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B1 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A1 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A2 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A3 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A5 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B2 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B2 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B4 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B5 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C2 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C6 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B6 = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D1 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D2 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D3 = CLBLM_L_X10Y117_SLICE_X13Y117_DQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D5 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A1 = CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A5 = CLBLM_L_X8Y117_SLICE_X11Y117_C5Q;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B1 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B6 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C3 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C1 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C5 = CLBLM_L_X10Y117_SLICE_X13Y117_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C6 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C6 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D1 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D2 = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D3 = CLBLM_R_X11Y119_SLICE_X14Y119_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D5 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D6 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A1 = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A2 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A4 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A5 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A6 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B2 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B3 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B4 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B5 = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B6 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C2 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C4 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D2 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D4 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A1 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A3 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A4 = CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A6 = CLBLM_L_X12Y119_SLICE_X16Y119_CQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B2 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B3 = CLBLM_R_X7Y114_SLICE_X9Y114_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B4 = CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B5 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B6 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C1 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C4 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C5 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C6 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D1 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D2 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D3 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D4 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D5 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D6 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X37Y120_SLICE_X56Y120_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A1 = CLBLM_L_X10Y117_SLICE_X13Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A3 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A4 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_AX = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B1 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B2 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B4 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C1 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C6 = CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D5 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D6 = CLBLM_R_X7Y116_SLICE_X9Y116_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A2 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A4 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A5 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B4 = CLBLM_R_X7Y116_SLICE_X9Y116_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C3 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C5 = CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D3 = CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D5 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A1 = CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A2 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A3 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A4 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A5 = CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A6 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C1 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C2 = CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C3 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C4 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C5 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C6 = CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D1 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D2 = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D3 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D4 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D5 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D6 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A1 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A2 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A3 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A5 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A6 = CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B1 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B2 = CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B3 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B5 = CLBLM_R_X13Y121_SLICE_X18Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C1 = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C2 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C3 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C4 = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C5 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C6 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D1 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D2 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D4 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D5 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D6 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = CLBLM_R_X11Y118_SLICE_X15Y118_DQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_DQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_B5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_AX = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = CLBLM_R_X11Y119_SLICE_X14Y119_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = CLBLM_R_X3Y119_SLICE_X2Y119_B5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A1 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A2 = CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A3 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B1 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B2 = CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B3 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B4 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B5 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B6 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C3 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C4 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D1 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D2 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D3 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D4 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D5 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A1 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A3 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A5 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B1 = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B2 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B4 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B5 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B6 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C1 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C2 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C3 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C4 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C5 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D1 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D2 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D3 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D4 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D5 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D6 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C2 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C4 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C5 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_AX = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = CLBLM_R_X11Y119_SLICE_X14Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = CLBLM_R_X5Y114_SLICE_X7Y114_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_SR = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = CLBLM_R_X5Y115_SLICE_X6Y115_DQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = CLBLM_R_X5Y115_SLICE_X6Y115_DQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A1 = CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A2 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A4 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A5 = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A6 = CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B2 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B3 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B4 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B5 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A3 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C1 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C2 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C3 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B1 = CLBLM_L_X8Y120_SLICE_X11Y120_DQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B2 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B3 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C4 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C5 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_B5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = CLBLM_L_X10Y123_SLICE_X12Y123_DQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B2 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D1 = CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D2 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D3 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_B5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_AX = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = CLBLM_L_X10Y118_SLICE_X12Y118_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_DX = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A2 = CLBLM_L_X12Y115_SLICE_X17Y115_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A3 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A5 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B2 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B6 = CLBLM_L_X12Y116_SLICE_X16Y116_CQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B6 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A1 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A2 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A4 = CLBLM_R_X5Y114_SLICE_X7Y114_DQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A5 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_AX = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B1 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B2 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B5 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C2 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C4 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C5 = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C6 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C6 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D1 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D2 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D3 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D4 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D5 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D6 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_AX = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A1 = CLBLM_L_X10Y122_SLICE_X12Y122_DQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A2 = CLBLM_L_X10Y120_SLICE_X13Y120_DQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A3 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A4 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B1 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B2 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B3 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B4 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B6 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B2 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C1 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C2 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C3 = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D3 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D4 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D5 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A2 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_A5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A5 = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B2 = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_D5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C3 = CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C4 = CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D2 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B2 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B5 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A2 = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A4 = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A5 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C4 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B1 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B3 = CLBLM_L_X12Y115_SLICE_X17Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B4 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B5 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B6 = CLBLM_L_X12Y116_SLICE_X16Y116_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C1 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C2 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C3 = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C4 = CLBLM_L_X12Y116_SLICE_X16Y116_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D2 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D3 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D5 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A1 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A3 = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A4 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A5 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B1 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B2 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B4 = CLBLM_L_X8Y113_SLICE_X11Y113_B5Q;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B5 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B6 = CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D2 = CLBLM_R_X11Y121_SLICE_X15Y121_CQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C1 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C4 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D3 = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D4 = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D5 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D2 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D3 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D4 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D6 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D6 = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_A3 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_A4 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_B2 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_B3 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_B5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A1 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A4 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A6 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C4 = CLBLM_R_X7Y123_SLICE_X8Y123_D5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B2 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B5 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C5 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C2 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C4 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D2 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D4 = CLBLM_L_X10Y117_SLICE_X13Y117_DQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A1 = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A2 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A3 = CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A4 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_AX = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B1 = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B3 = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B4 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B5 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C3 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C4 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D1 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D5 = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_A5Q;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A1 = CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A2 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A4 = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A6 = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B4 = CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B5 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_C6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C2 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C3 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C5 = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D1 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D2 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D3 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C5 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D6 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A5 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A6 = CLBLM_L_X12Y116_SLICE_X16Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B1 = CLBLM_L_X10Y118_SLICE_X13Y118_DQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B5 = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B6 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C1 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C3 = CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C5 = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D4 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D2 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D3 = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D4 = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D6 = 1'b1;
  assign CLBLM_R_X37Y120_SLICE_X57Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D2 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D3 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C5 = CLBLM_R_X7Y123_SLICE_X9Y123_DQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D3 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_DQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = CLBLM_R_X7Y123_SLICE_X9Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_AX = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = CLBLM_L_X8Y120_SLICE_X11Y120_DQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_A5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = CLBLM_L_X8Y123_SLICE_X10Y123_D5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = CLBLL_L_X4Y118_SLICE_X4Y118_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = CLBLM_R_X7Y116_SLICE_X9Y116_CQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = CLBLM_R_X7Y114_SLICE_X9Y114_B5Q;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = CLBLM_R_X5Y120_SLICE_X7Y120_B5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = CLBLL_L_X4Y118_SLICE_X4Y118_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = CLBLL_L_X4Y118_SLICE_X4Y118_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A2 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A4 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B2 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B4 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B6 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C5 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C1 = CLBLM_R_X11Y117_SLICE_X15Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C2 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C4 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D1 = CLBLM_R_X7Y116_SLICE_X9Y116_CQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D3 = CLBLM_R_X11Y117_SLICE_X15Y117_DQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D4 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A2 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A3 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B1 = CLBLM_R_X11Y121_SLICE_X15Y121_CQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B2 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B4 = CLBLM_L_X10Y120_SLICE_X12Y120_D5Q;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C2 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C4 = CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C5 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D2 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_C5Q;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D4 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_DQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A1 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A2 = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A3 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A4 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A5 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A6 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B1 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B4 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B6 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = CLBLM_R_X5Y113_SLICE_X7Y113_B5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C1 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C2 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C3 = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C6 = CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D3 = CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D4 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D5 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A3 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A6 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B4 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = CLBLM_R_X3Y116_SLICE_X2Y116_CQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C4 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D1 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D3 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D4 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D5 = CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D6 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = CLBLM_R_X5Y114_SLICE_X7Y114_DQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = CLBLM_L_X12Y116_SLICE_X16Y116_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A5 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A6 = CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B1 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B2 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B4 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B5 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C2 = CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C3 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C4 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C5 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D3 = CLBLM_R_X11Y118_SLICE_X15Y118_DQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D4 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D5 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D6 = CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A1 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A2 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A3 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A4 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A5 = CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B1 = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B2 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B4 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B5 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B6 = CLBLM_R_X3Y117_SLICE_X3Y117_CQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C1 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C4 = CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D1 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D2 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D3 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D4 = CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D5 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_D5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C4 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B1 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B2 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B3 = CLBLM_L_X8Y117_SLICE_X11Y117_DQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A2 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A3 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A4 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A5 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B1 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B2 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B3 = CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B5 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A1 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A2 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C1 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C4 = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C5 = CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C6 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C1 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A4 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A6 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D1 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C6 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D2 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D3 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C3 = CLBLM_L_X8Y113_SLICE_X11Y113_B5Q;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D2 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C6 = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A1 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A2 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A4 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A5 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D2 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D3 = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D4 = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D5 = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D6 = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B4 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B5 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_C5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D5 = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C5 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A5 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B6 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D2 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D4 = CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D5 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D6 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C5 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_SR = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B1 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B2 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B3 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B6 = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D4 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D6 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D5 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A5 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A1 = CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A2 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A4 = CLBLM_L_X12Y117_SLICE_X16Y117_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A6 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B1 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C1 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C4 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D1 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D3 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D4 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A2 = CLBLM_R_X11Y119_SLICE_X14Y119_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A3 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A5 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B2 = CLBLM_R_X11Y119_SLICE_X14Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B4 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C4 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C6 = CLBLM_R_X13Y122_SLICE_X18Y122_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D1 = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D3 = CLBLM_R_X11Y119_SLICE_X14Y119_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D5 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D1 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A4 = CLBLM_L_X12Y121_SLICE_X17Y121_BQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D4 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A1 = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A2 = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A3 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A4 = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A5 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A6 = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A5 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B1 = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B2 = CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B4 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C1 = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B6 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C6 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_B5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = CLBLM_R_X7Y116_SLICE_X9Y116_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D4 = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D5 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A4 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A5 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B5 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C1 = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C4 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C6 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C5 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = CLBLM_R_X11Y119_SLICE_X14Y119_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = CLBLM_R_X7Y122_SLICE_X9Y122_DQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D1 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D2 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D3 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D4 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A1 = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A3 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A4 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A6 = CLBLM_R_X11Y121_SLICE_X15Y121_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C2 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C3 = CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B1 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B2 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B3 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B4 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B6 = CLBLM_R_X5Y115_SLICE_X6Y115_DQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C4 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C5 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C4 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C5 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C6 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C6 = CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D2 = CLBLM_L_X12Y120_SLICE_X16Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D4 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D5 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D6 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A1 = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A3 = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A5 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B1 = CLBLM_R_X11Y120_SLICE_X15Y120_DQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B2 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B3 = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C1 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C2 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C3 = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D1 = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D1 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D3 = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D6 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D5 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A1 = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A2 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A3 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A6 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B1 = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B3 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B4 = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B5 = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B6 = CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C4 = CLBLL_L_X2Y119_SLICE_X1Y119_A5Q;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A2 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A3 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C4 = CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A4 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C5 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B1 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B2 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D4 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D2 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C2 = CLBLM_L_X8Y117_SLICE_X11Y117_CQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C5 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B5 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B6 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D1 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D2 = CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D3 = CLBLM_L_X8Y117_SLICE_X11Y117_DQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D4 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D6 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A2 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A4 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A1 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A2 = CLBLM_R_X7Y123_SLICE_X9Y123_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A4 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A5 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B5 = CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B6 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C1 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C3 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D2 = CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D5 = CLBLM_R_X7Y119_SLICE_X8Y119_B5Q;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D1 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D2 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D3 = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D4 = CLBLM_L_X8Y117_SLICE_X11Y117_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D5 = CLBLM_L_X10Y117_SLICE_X12Y117_DQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D6 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A2 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A4 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B1 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B4 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B6 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B2 = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B3 = CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C5 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C6 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B4 = CLBLM_L_X12Y120_SLICE_X16Y120_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D1 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A3 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A4 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A1 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_AX = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B1 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B2 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B6 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C2 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B5 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C4 = CLBLM_R_X11Y121_SLICE_X14Y121_A5Q;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C6 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B6 = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D2 = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D4 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D5 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D6 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C4 = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C5 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A2 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B1 = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B2 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A1 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A3 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A4 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A6 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_A5Q;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B5 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B6 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C2 = CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C4 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A2 = CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D3 = CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D4 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D6 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A2 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A4 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A5 = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A4 = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B3 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B5 = CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B1 = CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C2 = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C3 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B2 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C5 = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C6 = CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D3 = CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B4 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D5 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D6 = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A1 = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A3 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B1 = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B2 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B3 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B5 = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C3 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = CLBLM_R_X7Y114_SLICE_X9Y114_DQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C4 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C5 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C6 = CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D3 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A6 = CLBLM_R_X11Y120_SLICE_X15Y120_DQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B1 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B3 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C1 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C2 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D1 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D2 = CLBLM_L_X8Y122_SLICE_X10Y122_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D3 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D6 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D4 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B4 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B5 = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B6 = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C4 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A3 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A4 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A5 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A6 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C6 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C1 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C2 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A2 = CLBLM_L_X10Y122_SLICE_X12Y122_A5Q;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B5 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_AX = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B3 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C3 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D2 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D3 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D5 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A1 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A2 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A4 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A5 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A6 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B1 = CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B2 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B3 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B4 = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B5 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B6 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D1 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D2 = CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = CLBLM_R_X7Y114_SLICE_X9Y114_DQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D3 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D4 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A1 = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A2 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A3 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A4 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A5 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B1 = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B3 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B4 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B5 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B6 = CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C1 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C2 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C3 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D1 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = CLBLM_R_X7Y114_SLICE_X9Y114_B5Q;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D2 = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D3 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D4 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D6 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_SR = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B6 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A3 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A4 = CLBLM_L_X10Y120_SLICE_X12Y120_C5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A6 = CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B4 = CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B2 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C1 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C2 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C5 = CLBLM_L_X10Y123_SLICE_X12Y123_D5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A2 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A4 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D3 = CLBLM_L_X8Y120_SLICE_X11Y120_DQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D4 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D6 = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A2 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A4 = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A6 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_AX = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B3 = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C2 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C4 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D1 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D3 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D5 = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A1 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A3 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A4 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B1 = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B4 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B6 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = CLBLM_R_X7Y114_SLICE_X9Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = CLBLM_R_X7Y123_SLICE_X8Y123_D5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C2 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C3 = CLBLM_R_X11Y124_SLICE_X15Y124_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_B5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D3 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D4 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A3 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A4 = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = CLBLM_R_X7Y114_SLICE_X9Y114_DQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = CLBLM_R_X11Y118_SLICE_X15Y118_DQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A6 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B1 = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B3 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B4 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C1 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C2 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_BX = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D2 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D3 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D4 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D5 = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D6 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B1 = CLBLM_R_X13Y120_SLICE_X18Y120_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B2 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_CX = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B3 = CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B4 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B5 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B6 = CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A2 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A4 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A5 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A6 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B1 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C2 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C5 = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D1 = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D4 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A3 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B2 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B3 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B4 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B5 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B6 = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C6 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D1 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D2 = CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D4 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D6 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A4 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = CLBLM_R_X7Y124_SLICE_X9Y124_DQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_AX = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A1 = CLBLM_L_X8Y117_SLICE_X11Y117_DQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A3 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A4 = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B3 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B4 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D4 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D5 = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D6 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X10Y123_SLICE_X12Y123_D5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A1 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A3 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A5 = CLBLM_L_X8Y121_SLICE_X11Y121_A5Q;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_AX = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B5 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B6 = CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C4 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C5 = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D1 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D3 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D4 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D5 = CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D6 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A3 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B2 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B4 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A6 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C1 = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C2 = CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C5 = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B2 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B3 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C2 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D2 = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D3 = CLBLM_L_X8Y122_SLICE_X10Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D6 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C5 = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C6 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = CLBLM_L_X8Y124_SLICE_X10Y124_D5Q;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = CLBLM_R_X7Y116_SLICE_X9Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D5 = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_B5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = CLBLM_R_X7Y116_SLICE_X8Y116_DQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = CLBLM_R_X7Y114_SLICE_X9Y114_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A5 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X4Y118_SLICE_X4Y118_CQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A1 = CLBLM_L_X8Y123_SLICE_X10Y123_DQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A3 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A4 = CLBLM_L_X10Y120_SLICE_X13Y120_DQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A5 = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B1 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B2 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B3 = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B4 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B5 = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B6 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C1 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C2 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C3 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C4 = CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C5 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C6 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D1 = CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A1 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A3 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A4 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B6 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C5 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C2 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D2 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D4 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = CLBLM_R_X7Y116_SLICE_X9Y116_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C3 = CLBLM_R_X3Y119_SLICE_X2Y119_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D1 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C5 = CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C6 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A4 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A5 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A6 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D3 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C4 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_AX = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B2 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B4 = CLBLM_R_X3Y116_SLICE_X2Y116_CQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B5 = CLBLM_L_X10Y122_SLICE_X13Y122_D5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C1 = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C2 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C3 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C4 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D2 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D3 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D4 = CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D4 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D4 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D5 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A1 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A2 = CLBLM_L_X10Y122_SLICE_X13Y122_D5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A4 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B2 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B3 = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B5 = CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C1 = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C2 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D2 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D5 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D6 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A3 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B1 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B5 = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B6 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C4 = CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C5 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C6 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D3 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D6 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A1 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A2 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A3 = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A5 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A6 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A3 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B1 = CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B5 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B6 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C1 = CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C2 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C3 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A6 = CLBLL_L_X4Y125_SLICE_X5Y125_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C6 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D1 = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D2 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D3 = CLBLM_L_X8Y118_SLICE_X11Y118_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D4 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D5 = CLBLM_L_X12Y119_SLICE_X16Y119_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B4 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B6 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A1 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A2 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A4 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A5 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B2 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B3 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B4 = CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B6 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C2 = CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C3 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C4 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C5 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D3 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D4 = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D5 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A1 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A4 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B1 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B5 = CLBLM_R_X5Y125_SLICE_X6Y125_DQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B6 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C1 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C2 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C3 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C5 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D1 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D3 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D5 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D6 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A1 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A4 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B2 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B3 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B4 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B5 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_AX = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D5 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A3 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A4 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A5 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = CLBLM_R_X7Y119_SLICE_X9Y119_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B2 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B3 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D6 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C3 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D1 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D5 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C4 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C6 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C2 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A4 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D6 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_DQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = CLBLM_R_X11Y121_SLICE_X14Y121_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C6 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = CLBLM_R_X7Y122_SLICE_X9Y122_DQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = CLBLM_R_X7Y119_SLICE_X9Y119_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = CLBLM_L_X12Y119_SLICE_X16Y119_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D2 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = CLBLM_R_X11Y121_SLICE_X14Y121_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D5 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D1 = CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D6 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D2 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D4 = CLBLM_L_X12Y122_SLICE_X17Y122_BQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = CLBLM_R_X7Y119_SLICE_X9Y119_A5Q;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B6 = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AX = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = CLBLM_R_X3Y120_SLICE_X3Y120_CQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = CLBLL_L_X2Y119_SLICE_X1Y119_A5Q;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C5 = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C6 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_AX = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B5 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B4 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B5 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_AX = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C4 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_AX = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A1 = CLBLM_L_X8Y120_SLICE_X11Y120_DQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A2 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B1 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A1 = CLBLM_L_X10Y124_SLICE_X12Y124_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A3 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A5 = CLBLM_R_X11Y119_SLICE_X14Y119_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B2 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B4 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B5 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B6 = CLBLM_L_X10Y122_SLICE_X12Y122_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C2 = CLBLM_R_X7Y123_SLICE_X9Y123_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C3 = CLBLM_L_X8Y122_SLICE_X11Y122_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_BX = CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D1 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D3 = CLBLM_R_X7Y123_SLICE_X9Y123_DQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D4 = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A1 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A2 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A4 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B1 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B2 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B3 = CLBLM_R_X7Y123_SLICE_X8Y123_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = CLBLM_R_X5Y124_SLICE_X7Y124_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C2 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D5 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C5 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A3 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A4 = CLBLM_R_X29Y141_SLICE_X42Y141_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A6 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A2 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B3 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = CLBLM_R_X11Y124_SLICE_X15Y124_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D3 = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D4 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D6 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_BX = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A1 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A3 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A5 = CLBLM_L_X10Y124_SLICE_X12Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B1 = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B2 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B4 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B6 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C2 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D2 = CLBLM_R_X7Y124_SLICE_X9Y124_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_C5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D3 = CLBLM_R_X7Y124_SLICE_X9Y124_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D4 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A2 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A5 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = CLBLM_R_X5Y114_SLICE_X7Y114_DQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = CLBLM_R_X7Y116_SLICE_X9Y116_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B1 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B4 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C1 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C2 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C3 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D2 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D3 = CLBLM_L_X8Y124_SLICE_X11Y124_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D4 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D5 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D6 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B4 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X8Y124_SLICE_X10Y124_DQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A4 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C4 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B3 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B6 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C1 = CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C2 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C3 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C4 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C5 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C6 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C6 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B5 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C2 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = CLBLL_L_X4Y118_SLICE_X4Y118_C5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D5 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C4 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C5 = CLBLM_L_X12Y123_SLICE_X16Y123_CQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = CLBLM_R_X5Y115_SLICE_X6Y115_DQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C6 = CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A3 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A4 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A6 = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B6 = CLBLM_R_X29Y141_SLICE_X42Y141_AO6;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C1 = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D1 = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D3 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A1 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B6 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A2 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A3 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B2 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B3 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A5 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C1 = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C2 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C3 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C4 = CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C5 = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C6 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A6 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D1 = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D2 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D3 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D4 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D5 = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D6 = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A1 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A3 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A4 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A4 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A5 = CLBLM_L_X8Y125_SLICE_X10Y125_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A6 = CLBLM_R_X7Y119_SLICE_X8Y119_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B1 = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = CLBLM_R_X11Y119_SLICE_X14Y119_DQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = CLBLM_R_X11Y117_SLICE_X15Y117_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A1 = CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = CLBLM_L_X10Y122_SLICE_X13Y122_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B2 = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B3 = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B5 = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B1 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y124_SLICE_X10Y124_D5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = CLBLL_L_X4Y118_SLICE_X5Y118_DQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = CLBLM_R_X7Y116_SLICE_X9Y116_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C4 = CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X5Y115_SLICE_X7Y115_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = CLBLM_R_X7Y123_SLICE_X8Y123_D5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X10Y123_SLICE_X12Y123_D5Q;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = CLBLM_R_X5Y114_SLICE_X7Y114_DQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = CLBLM_L_X8Y121_SLICE_X11Y121_B5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = CLBLM_R_X7Y123_SLICE_X8Y123_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = CLBLM_R_X7Y123_SLICE_X8Y123_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = CLBLM_R_X7Y123_SLICE_X8Y123_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_AX = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = CLBLL_L_X4Y118_SLICE_X5Y118_DQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_DQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = CLBLM_R_X7Y122_SLICE_X9Y122_DQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = CLBLM_R_X3Y116_SLICE_X2Y116_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = CLBLM_R_X11Y121_SLICE_X14Y121_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = CLBLM_R_X5Y113_SLICE_X7Y113_B5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A3 = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A4 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B1 = CLBLM_R_X11Y121_SLICE_X15Y121_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B2 = CLBLM_R_X5Y121_SLICE_X7Y121_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B3 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B5 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B6 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C2 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C3 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C4 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C5 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D4 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D5 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A2 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A4 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B1 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B2 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C1 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C4 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C5 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D1 = CLBLM_R_X29Y141_SLICE_X42Y141_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D2 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D3 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D6 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_BX = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D2 = CLBLM_L_X10Y120_SLICE_X13Y120_DQ;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A1 = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A3 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = CLBLM_L_X12Y119_SLICE_X16Y119_BQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y115_SLICE_X18Y115_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A1 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A3 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A4 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A6 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C1 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B2 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B3 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B4 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B6 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C2 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C3 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C4 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C6 = CLBLM_L_X8Y123_SLICE_X10Y123_D5Q;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D2 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D3 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D5 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D6 = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A1 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A3 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A4 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A6 = CLBLM_R_X5Y125_SLICE_X6Y125_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B1 = CLBLM_L_X10Y122_SLICE_X12Y122_B5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B5 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B6 = CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C1 = CLBLM_R_X29Y141_SLICE_X42Y141_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C3 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C4 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C6 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D1 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D3 = CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D4 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D6 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A1 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A2 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A6 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B2 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B4 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C2 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C6 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D2 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D5 = CLBLM_R_X7Y124_SLICE_X9Y124_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D6 = CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A3 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B1 = CLBLM_R_X7Y123_SLICE_X9Y123_DQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B2 = CLBLM_R_X29Y141_SLICE_X42Y141_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B4 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C1 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C4 = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C6 = CLBLM_R_X29Y141_SLICE_X42Y141_AO6;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D3 = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D4 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D5 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D6 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A4 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B2 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B4 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C2 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C4 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C6 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D3 = CLBLM_R_X5Y124_SLICE_X7Y124_DQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D5 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D6 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A1 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A2 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A4 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A5 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A6 = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B1 = CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B2 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B3 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B5 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B6 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_BX = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C1 = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C2 = CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C4 = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C5 = CLBLM_R_X5Y124_SLICE_X7Y124_DQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C6 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = CLBLL_L_X2Y119_SLICE_X1Y119_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_BX = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X37Y120_SLICE_X56Y120_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A5 = CLBLM_L_X8Y117_SLICE_X11Y117_C5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = CLBLM_L_X10Y118_SLICE_X12Y118_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C1 = CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_A1 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_A2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_A6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_B1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_B4 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_D5Q;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_B6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_C1 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_C2 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_C3 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_C4 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_C5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_D1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_D2 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_D3 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_D5 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X43Y141_D6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C3 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_A3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_A4 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_A6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_B1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_B2 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_B3 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_B4 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_B5 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_B6 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_C1 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_C2 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_C3 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_C4 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_C5 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_C6 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_D1 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_D2 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_D3 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_D4 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_D5 = 1'b1;
  assign CLBLM_R_X29Y141_SLICE_X42Y141_D6 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A1 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A2 = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A6 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B1 = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B2 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B4 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B5 = CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AX = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C3 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_L_X12Y116_SLICE_X16Y116_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLM_R_X5Y115_SLICE_X6Y115_DQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A2 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A6 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B1 = CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D1 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D2 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D3 = CLBLM_R_X5Y125_SLICE_X6Y125_DQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D6 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = 1'b1;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D1 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D2 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AX = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = CLBLM_R_X7Y124_SLICE_X9Y124_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = CLBLM_R_X3Y116_SLICE_X2Y116_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = CLBLM_R_X5Y113_SLICE_X7Y113_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = CLBLM_R_X3Y121_SLICE_X3Y121_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = CLBLM_R_X5Y113_SLICE_X7Y113_B5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D5 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D6 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X29Y141_SLICE_X42Y141_AO5;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X29Y141_SLICE_X42Y141_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B2 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B3 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B4 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = CLBLM_R_X3Y117_SLICE_X3Y117_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = CLBLM_R_X3Y117_SLICE_X2Y117_CQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = CLBLM_R_X3Y116_SLICE_X2Y116_C5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = CLBLL_L_X4Y116_SLICE_X4Y116_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = CLBLM_R_X3Y117_SLICE_X2Y117_DQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = CLBLM_L_X8Y120_SLICE_X10Y120_C5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = CLBLM_L_X8Y114_SLICE_X11Y114_A5Q;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLM_R_X7Y116_SLICE_X8Y116_DQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = CLBLL_L_X4Y119_SLICE_X4Y119_A5Q;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = CLBLL_L_X2Y119_SLICE_X1Y119_A5Q;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = CLBLM_L_X8Y114_SLICE_X11Y114_A5Q;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = CLBLM_L_X8Y113_SLICE_X11Y113_DQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = CLBLM_L_X10Y116_SLICE_X13Y116_A5Q;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C4 = 1'b1;
endmodule
