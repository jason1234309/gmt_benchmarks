module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_SING_X0Y149_IOB_X0Y149_IPAD,
  input LIOB33_SING_X0Y150_IOB_X0Y150_IPAD,
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_SING_X0Y99_IOB_X0Y99_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input LIOB33_X0Y123_IOB_X0Y124_IPAD,
  input LIOB33_X0Y125_IOB_X0Y125_IPAD,
  input LIOB33_X0Y125_IOB_X0Y126_IPAD,
  input LIOB33_X0Y127_IOB_X0Y127_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  input LIOB33_X0Y129_IOB_X0Y129_IPAD,
  input LIOB33_X0Y129_IOB_X0Y130_IPAD,
  input LIOB33_X0Y131_IOB_X0Y131_IPAD,
  input LIOB33_X0Y131_IOB_X0Y132_IPAD,
  input LIOB33_X0Y133_IOB_X0Y133_IPAD,
  input LIOB33_X0Y133_IOB_X0Y134_IPAD,
  input LIOB33_X0Y135_IOB_X0Y135_IPAD,
  input LIOB33_X0Y135_IOB_X0Y136_IPAD,
  input LIOB33_X0Y137_IOB_X0Y137_IPAD,
  input LIOB33_X0Y137_IOB_X0Y138_IPAD,
  input LIOB33_X0Y139_IOB_X0Y139_IPAD,
  input LIOB33_X0Y139_IOB_X0Y140_IPAD,
  input LIOB33_X0Y141_IOB_X0Y141_IPAD,
  input LIOB33_X0Y141_IOB_X0Y142_IPAD,
  input LIOB33_X0Y143_IOB_X0Y143_IPAD,
  input LIOB33_X0Y145_IOB_X0Y145_IPAD,
  input LIOB33_X0Y145_IOB_X0Y146_IPAD,
  input LIOB33_X0Y147_IOB_X0Y147_IPAD,
  input LIOB33_X0Y147_IOB_X0Y148_IPAD,
  input LIOB33_X0Y151_IOB_X0Y151_IPAD,
  input LIOB33_X0Y151_IOB_X0Y152_IPAD,
  input LIOB33_X0Y153_IOB_X0Y153_IPAD,
  input LIOB33_X0Y153_IOB_X0Y154_IPAD,
  input LIOB33_X0Y155_IOB_X0Y155_IPAD,
  input LIOB33_X0Y155_IOB_X0Y156_IPAD,
  input LIOB33_X0Y157_IOB_X0Y157_IPAD,
  input LIOB33_X0Y157_IOB_X0Y158_IPAD,
  input LIOB33_X0Y159_IOB_X0Y159_IPAD,
  input LIOB33_X0Y159_IOB_X0Y160_IPAD,
  input LIOB33_X0Y161_IOB_X0Y161_IPAD,
  input LIOB33_X0Y161_IOB_X0Y162_IPAD,
  input LIOB33_X0Y163_IOB_X0Y163_IPAD,
  input LIOB33_X0Y163_IOB_X0Y164_IPAD,
  input LIOB33_X0Y165_IOB_X0Y165_IPAD,
  input LIOB33_X0Y165_IOB_X0Y166_IPAD,
  input LIOB33_X0Y167_IOB_X0Y167_IPAD,
  input LIOB33_X0Y167_IOB_X0Y168_IPAD,
  input LIOB33_X0Y169_IOB_X0Y169_IPAD,
  input LIOB33_X0Y169_IOB_X0Y170_IPAD,
  input LIOB33_X0Y171_IOB_X0Y171_IPAD,
  input LIOB33_X0Y171_IOB_X0Y172_IPAD,
  input LIOB33_X0Y173_IOB_X0Y173_IPAD,
  input LIOB33_X0Y173_IOB_X0Y174_IPAD,
  input LIOB33_X0Y175_IOB_X0Y175_IPAD,
  input LIOB33_X0Y175_IOB_X0Y176_IPAD,
  input LIOB33_X0Y177_IOB_X0Y177_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input LIOB33_X0Y79_IOB_X0Y80_IPAD,
  input LIOB33_X0Y81_IOB_X0Y81_IPAD,
  input LIOB33_X0Y81_IOB_X0Y82_IPAD,
  input LIOB33_X0Y83_IOB_X0Y83_IPAD,
  input LIOB33_X0Y83_IOB_X0Y84_IPAD,
  input LIOB33_X0Y85_IOB_X0Y85_IPAD,
  input LIOB33_X0Y85_IOB_X0Y86_IPAD,
  input LIOB33_X0Y87_IOB_X0Y87_IPAD,
  input LIOB33_X0Y87_IOB_X0Y88_IPAD,
  input LIOB33_X0Y89_IOB_X0Y89_IPAD,
  input LIOB33_X0Y89_IOB_X0Y90_IPAD,
  input LIOB33_X0Y91_IOB_X0Y91_IPAD,
  input LIOB33_X0Y91_IOB_X0Y92_IPAD,
  input LIOB33_X0Y93_IOB_X0Y93_IPAD,
  input LIOB33_X0Y93_IOB_X0Y94_IPAD,
  input LIOB33_X0Y95_IOB_X0Y95_IPAD,
  input LIOB33_X0Y95_IOB_X0Y96_IPAD,
  input LIOB33_X0Y97_IOB_X0Y97_IPAD,
  input LIOB33_X0Y97_IOB_X0Y98_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y150_IOB_X1Y150_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y151_IOB_X1Y151_IPAD,
  input RIOB33_X105Y151_IOB_X1Y152_IPAD,
  input RIOB33_X105Y153_IOB_X1Y153_IPAD,
  input RIOB33_X105Y153_IOB_X1Y154_IPAD,
  input RIOB33_X105Y155_IOB_X1Y155_IPAD,
  input RIOB33_X105Y155_IOB_X1Y156_IPAD,
  input RIOB33_X105Y157_IOB_X1Y157_IPAD,
  input RIOB33_X105Y157_IOB_X1Y158_IPAD,
  input RIOB33_X105Y159_IOB_X1Y159_IPAD,
  input RIOB33_X105Y159_IOB_X1Y160_IPAD,
  input RIOB33_X105Y161_IOB_X1Y161_IPAD,
  input RIOB33_X105Y161_IOB_X1Y162_IPAD,
  input RIOB33_X105Y163_IOB_X1Y163_IPAD,
  input RIOB33_X105Y163_IOB_X1Y164_IPAD,
  input RIOB33_X105Y165_IOB_X1Y165_IPAD,
  input RIOB33_X105Y165_IOB_X1Y166_IPAD,
  input RIOB33_X105Y167_IOB_X1Y167_IPAD,
  input RIOB33_X105Y167_IOB_X1Y168_IPAD,
  input RIOB33_X105Y169_IOB_X1Y169_IPAD,
  input RIOB33_X105Y169_IOB_X1Y170_IPAD,
  input RIOB33_X105Y171_IOB_X1Y171_IPAD,
  input RIOB33_X105Y171_IOB_X1Y172_IPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_SING_X0Y200_IOB_X0Y200_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output RIOB33_SING_X105Y149_IOB_X1Y149_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_SING_X105Y50_IOB_X1Y50_OPAD,
  output RIOB33_SING_X105Y99_IOB_X1Y99_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y127_IOB_X1Y128_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD,
  output RIOB33_X105Y145_IOB_X1Y146_OPAD,
  output RIOB33_X105Y147_IOB_X1Y147_OPAD,
  output RIOB33_X105Y147_IOB_X1Y148_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD,
  output RIOB33_X105Y51_IOB_X1Y51_OPAD,
  output RIOB33_X105Y51_IOB_X1Y52_OPAD,
  output RIOB33_X105Y53_IOB_X1Y53_OPAD,
  output RIOB33_X105Y53_IOB_X1Y54_OPAD,
  output RIOB33_X105Y55_IOB_X1Y55_OPAD,
  output RIOB33_X105Y55_IOB_X1Y56_OPAD,
  output RIOB33_X105Y57_IOB_X1Y57_OPAD,
  output RIOB33_X105Y57_IOB_X1Y58_OPAD,
  output RIOB33_X105Y59_IOB_X1Y59_OPAD,
  output RIOB33_X105Y59_IOB_X1Y60_OPAD,
  output RIOB33_X105Y61_IOB_X1Y61_OPAD,
  output RIOB33_X105Y61_IOB_X1Y62_OPAD,
  output RIOB33_X105Y63_IOB_X1Y63_OPAD,
  output RIOB33_X105Y63_IOB_X1Y64_OPAD,
  output RIOB33_X105Y65_IOB_X1Y65_OPAD,
  output RIOB33_X105Y65_IOB_X1Y66_OPAD,
  output RIOB33_X105Y67_IOB_X1Y67_OPAD,
  output RIOB33_X105Y67_IOB_X1Y68_OPAD,
  output RIOB33_X105Y69_IOB_X1Y69_OPAD,
  output RIOB33_X105Y69_IOB_X1Y70_OPAD,
  output RIOB33_X105Y71_IOB_X1Y71_OPAD,
  output RIOB33_X105Y71_IOB_X1Y72_OPAD,
  output RIOB33_X105Y73_IOB_X1Y73_OPAD,
  output RIOB33_X105Y73_IOB_X1Y74_OPAD,
  output RIOB33_X105Y75_IOB_X1Y75_OPAD,
  output RIOB33_X105Y75_IOB_X1Y76_OPAD,
  output RIOB33_X105Y77_IOB_X1Y77_OPAD,
  output RIOB33_X105Y77_IOB_X1Y78_OPAD,
  output RIOB33_X105Y79_IOB_X1Y79_OPAD,
  output RIOB33_X105Y79_IOB_X1Y80_OPAD,
  output RIOB33_X105Y81_IOB_X1Y81_OPAD,
  output RIOB33_X105Y81_IOB_X1Y82_OPAD,
  output RIOB33_X105Y83_IOB_X1Y83_OPAD,
  output RIOB33_X105Y83_IOB_X1Y84_OPAD,
  output RIOB33_X105Y85_IOB_X1Y85_OPAD,
  output RIOB33_X105Y85_IOB_X1Y86_OPAD,
  output RIOB33_X105Y87_IOB_X1Y87_OPAD,
  output RIOB33_X105Y87_IOB_X1Y88_OPAD,
  output RIOB33_X105Y89_IOB_X1Y89_OPAD,
  output RIOB33_X105Y89_IOB_X1Y90_OPAD,
  output RIOB33_X105Y91_IOB_X1Y91_OPAD,
  output RIOB33_X105Y91_IOB_X1Y92_OPAD,
  output RIOB33_X105Y93_IOB_X1Y93_OPAD,
  output RIOB33_X105Y93_IOB_X1Y94_OPAD,
  output RIOB33_X105Y95_IOB_X1Y95_OPAD,
  output RIOB33_X105Y95_IOB_X1Y96_OPAD,
  output RIOB33_X105Y97_IOB_X1Y97_OPAD,
  output RIOB33_X105Y97_IOB_X1Y98_OPAD
  );
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_AO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_AO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_BO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_BO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_CO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_CO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_DO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_DO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_AO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_AO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_BO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_BO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_CO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_CO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_DO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_DO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A1;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A2;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A3;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A4;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_AO5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_AO6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A_CY;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_A_XOR;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B1;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B2;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B3;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B4;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_BO5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_BO6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B_CY;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_B_XOR;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C1;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C2;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C3;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C4;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_CO5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_CO6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C_CY;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_C_XOR;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D1;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D2;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D3;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D4;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_DO5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_DO6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D_CY;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X0Y101_D_XOR;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A1;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A2;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A3;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A4;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_AO5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_AO6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A_CY;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_A_XOR;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B1;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B2;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B3;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B4;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_BO5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_BO6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B_CY;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_B_XOR;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C1;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C2;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C3;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C4;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_CO5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_CO6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C_CY;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_C_XOR;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D1;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D2;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D3;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D4;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_DO5;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_DO6;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D_CY;
  wire [0:0] CLBLL_L_X2Y101_SLICE_X1Y101_D_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_AO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_AO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_BO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_CO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_CO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_DO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_DO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_AO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_AO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_BO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_BO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_CO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_CO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_DO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_DO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AMUX;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_AO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_BO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_BO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_CO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_CO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_DO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_DO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_AO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_BO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_CO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_CO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_DO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_DO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D_XOR;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A1;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A2;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A3;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A4;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_AMUX;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_AO5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_AO6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A_CY;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_A_XOR;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B1;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B2;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B3;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B4;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_BMUX;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_BO5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B_CY;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_B_XOR;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C1;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C2;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C3;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C4;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_CO5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_CO6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C_CY;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_C_XOR;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D1;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D2;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D3;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D4;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_DO5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_DO6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D_CY;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X0Y174_D_XOR;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A1;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A2;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A3;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A4;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_AO5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_AO6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A_CY;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_A_XOR;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B1;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B2;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B3;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B4;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_BO5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_BO6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B_CY;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_B_XOR;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C1;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C2;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C3;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C4;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_CO5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_CO6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C_CY;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_C_XOR;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D1;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D2;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D3;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D4;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_DO5;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_DO6;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D_CY;
  wire [0:0] CLBLL_L_X2Y174_SLICE_X1Y174_D_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_AO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_BO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_BO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_CO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_CO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_DO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_DO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_AO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_AO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_BO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_BO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_CO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_CO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_DO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_DO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D_XOR;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A1;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A2;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A3;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A4;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_AO5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_AO6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A_CY;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_A_XOR;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B1;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B2;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B3;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B4;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_BO5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_BO6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B_CY;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_B_XOR;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C1;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C2;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C3;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C4;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_CO5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_CO6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C_CY;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_C_XOR;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D1;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D2;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D3;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D4;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_DO5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_DO6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D_CY;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X126Y111_D_XOR;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A1;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A2;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A3;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A4;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_AO5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_AO6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A_CY;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_A_XOR;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B1;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B2;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B3;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B4;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_BO5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_BO6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B_CY;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_B_XOR;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C1;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C2;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C3;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C4;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_CO5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_CO6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C_CY;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_C_XOR;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D1;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D2;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D3;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D4;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_DO5;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_DO6;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D_CY;
  wire [0:0] CLBLL_R_X81Y111_SLICE_X127Y111_D_XOR;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A1;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A2;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A3;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A4;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_AO5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_AO6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A_CY;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_A_XOR;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B1;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B2;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B3;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B4;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_BO5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_BO6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B_CY;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_B_XOR;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C1;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C2;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C3;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C4;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_CO5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_CO6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C_CY;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_C_XOR;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D1;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D2;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D3;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D4;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_DO5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_DO6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D_CY;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X126Y122_D_XOR;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A1;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A2;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A3;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A4;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_AO5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_AO6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A_CY;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_A_XOR;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B1;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B2;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B3;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B4;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_BO5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_BO6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B_CY;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_B_XOR;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C1;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C2;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C3;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C4;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_CO5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_CO6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C_CY;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_C_XOR;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D1;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D2;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D3;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D4;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_DO5;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_DO6;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D_CY;
  wire [0:0] CLBLL_R_X81Y122_SLICE_X127Y122_D_XOR;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A1;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A2;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A3;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A4;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_AO5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_AO6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A_CY;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_A_XOR;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B1;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B2;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B3;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B4;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_BO5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_BO6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B_CY;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_B_XOR;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C1;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C2;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C3;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C4;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_CO5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_CO6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C_CY;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_C_XOR;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D1;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D2;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D3;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D4;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_DO5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_DO6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D_CY;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X126Y124_D_XOR;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A1;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A2;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A3;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A4;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_AO5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_AO6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A_CY;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_A_XOR;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B1;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B2;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B3;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B4;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_BO5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_BO6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B_CY;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_B_XOR;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C1;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C2;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C3;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C4;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_CO5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_CO6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C_CY;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_C_XOR;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D1;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D2;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D3;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D4;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_DO5;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_DO6;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D_CY;
  wire [0:0] CLBLL_R_X81Y124_SLICE_X127Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_XOR;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A1;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A2;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A3;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A4;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_AO5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_AO6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A_CY;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_A_XOR;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B1;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B2;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B3;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B4;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_BO5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_BO6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B_CY;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_B_XOR;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C1;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C2;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C3;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C4;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_CO5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_CO6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C_CY;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_C_XOR;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D1;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D2;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D3;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D4;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_DO5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_DO6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D_CY;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X44Y111_D_XOR;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A1;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A2;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A3;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A4;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_AO5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_AO6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A_CY;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_A_XOR;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B1;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B2;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B3;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B4;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_BO5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_BO6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B_CY;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_B_XOR;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C1;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C2;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C3;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C4;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_CO5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_CO6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C_CY;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_C_XOR;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D1;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D2;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D3;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D4;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_DO5;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_DO6;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D_CY;
  wire [0:0] CLBLM_L_X30Y111_SLICE_X45Y111_D_XOR;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A1;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A2;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A3;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A4;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_AO5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_AO6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A_CY;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_A_XOR;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B1;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B2;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B3;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B4;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_BO5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_BO6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B_CY;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_B_XOR;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C1;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C2;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C3;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C4;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_CO5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_CO6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C_CY;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_C_XOR;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D1;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D2;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D3;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D4;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_DO5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_DO6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D_CY;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X70Y121_D_XOR;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A1;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A2;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A3;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A4;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_AO5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_AO6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A_CY;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_A_XOR;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B1;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B2;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B3;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B4;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_BO5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_BO6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B_CY;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_B_XOR;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C1;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C2;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C3;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C4;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_CO5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_CO6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C_CY;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_C_XOR;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D1;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D2;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D3;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D4;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_DO5;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_DO6;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D_CY;
  wire [0:0] CLBLM_L_X46Y121_SLICE_X71Y121_D_XOR;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A1;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A2;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A3;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A4;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_AO5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_AO6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A_CY;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_A_XOR;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B1;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B2;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B3;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B4;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_BO5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_BO6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B_CY;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_B_XOR;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C1;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C2;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C3;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C4;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_CO5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_CO6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C_CY;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_C_XOR;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D1;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D2;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D3;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D4;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_DO5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_DO6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D_CY;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X70Y142_D_XOR;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A1;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A2;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A3;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A4;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_AO5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_AO6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A_CY;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_A_XOR;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B1;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B2;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B3;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B4;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_BO5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_BO6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B_CY;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_B_XOR;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C1;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C2;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C3;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C4;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_CO5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_CO6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C_CY;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_C_XOR;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D1;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D2;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D3;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D4;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_DO5;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_DO6;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D_CY;
  wire [0:0] CLBLM_L_X46Y142_SLICE_X71Y142_D_XOR;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A1;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A2;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A3;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A4;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_AMUX;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_AO5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_AO6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A_CY;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_A_XOR;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B1;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B2;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B3;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B4;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_BO5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_BO6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B_CY;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_B_XOR;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C1;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C2;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C3;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C4;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_CO5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_CO6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C_CY;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_C_XOR;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D1;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D2;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D3;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D4;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_DO5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_DO6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D_CY;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X76Y119_D_XOR;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A1;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A2;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A3;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A4;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_AO5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_AO6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A_CY;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_A_XOR;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B1;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B2;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B3;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B4;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_BO5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_BO6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B_CY;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_B_XOR;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C1;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C2;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C3;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C4;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_CO5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_CO6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C_CY;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_C_XOR;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D1;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D2;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D3;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D4;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_DO5;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_DO6;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D_CY;
  wire [0:0] CLBLM_L_X50Y119_SLICE_X77Y119_D_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_AO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_BO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_CO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_DO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_DO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_AO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_AO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_BO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_BO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_CO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_CO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_DO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_DO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D_XOR;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A1;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A2;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A3;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A4;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_AO5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_AO6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A_CY;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_A_XOR;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B1;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B2;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B3;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B4;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_BO5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_BO6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B_CY;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_B_XOR;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C1;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C2;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C3;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C4;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_CO5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_CO6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C_CY;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_C_XOR;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D1;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D2;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D3;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D4;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_DO5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_DO6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D_CY;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X120Y125_D_XOR;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A1;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A2;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A3;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A4;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_AO5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_AO6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A_CY;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_A_XOR;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B1;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B2;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B3;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B4;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_BO5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_BO6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B_CY;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_B_XOR;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C1;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C2;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C3;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C4;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_CO5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_CO6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C_CY;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_C_XOR;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D1;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D2;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D3;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D4;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_DO5;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_DO6;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D_CY;
  wire [0:0] CLBLM_L_X78Y125_SLICE_X121Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_AMUX;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_AO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_BMUX;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_BO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_CO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_CO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_DO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_DO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_AO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_AO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_BO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_BO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_CO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_CO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_DO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_DO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_AO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_AO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_BO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_BO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_CO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_CO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_DO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_DO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_AO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_AO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_BO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_BO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_CO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_CO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_DO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_DO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AMUX;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_BO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_CO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_DO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_AO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_BO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_DO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_DO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_AO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_AO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_BO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_BO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_CO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_DO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_AO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_AO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_BO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_BO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_CO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_CO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_DO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_DO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D_XOR;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A1;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A2;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A3;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A4;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_AO5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_AO6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A_CY;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_A_XOR;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B1;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B2;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B3;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B4;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_BO5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_BO6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B_CY;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_B_XOR;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C1;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C2;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C3;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C4;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_CO5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_CO6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C_CY;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_C_XOR;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D1;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D2;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D3;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D4;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_DO5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_DO6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D_CY;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X162Y103_D_XOR;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A1;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A2;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A3;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A4;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_AO5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_AO6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A_CY;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_A_XOR;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B1;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B2;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B3;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B4;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_BO5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_BO6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B_CY;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_B_XOR;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C1;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C2;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C3;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C4;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_CO5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_CO6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C_CY;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_C_XOR;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D1;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D2;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D3;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D4;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_DO5;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_DO6;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D_CY;
  wire [0:0] CLBLM_R_X103Y103_SLICE_X163Y103_D_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_AO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_AO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_BO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_BO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_CO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_CO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_DO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_DO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_AMUX;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_BO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_CO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_CO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_DO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_DO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_AO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_AO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_BO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_BO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_CO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_DO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_DO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AMUX;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_BO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_CO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_DO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_DO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_DO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_AO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_AO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_BO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_BO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_CO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_CO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_DO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_DO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_AMUX;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_AO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_AO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_BO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_BO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_CO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_CO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_DO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_DO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_AO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_AO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_BO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_BO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_CO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_CO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_DO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_DO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_AMUX;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_BO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_BO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_CO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_CO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_DO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_DO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_AO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_AO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_BO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_BO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_CO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_CO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_DO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_DO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_AO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_BO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_BO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_CO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_CO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_DO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_DO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_AO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_AO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_BO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_BO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_CO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_CO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_DO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_DO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_AO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_BO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_CO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_CO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_DO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_DO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_DO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_DO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AMUX;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BMUX;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_DO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_DO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_AO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_AO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_BO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_DO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_AMUX;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_AO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_BO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_BO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_CO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_CO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_DO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_DO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AMUX;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_DO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_DO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_DO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AMUX;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BMUX;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_DO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_AMUX;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_AO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_BO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_BO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_CO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_CO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_DO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_DO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_AO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_AO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_BO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_BO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_CO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_CO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_DO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_DO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_AMUX;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_AO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_AO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_BO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_CO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_CO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_DO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_DO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_AO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_AO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_BO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_BO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_CO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_CO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_DO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_DO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_AMUX;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_AO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_AO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_BO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_CO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_CO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_DO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_DO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_AMUX;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_AO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_AO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_BMUX;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_BO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_CO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_DO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_AO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_AO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_BO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_CO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_CO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_DO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_DO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_AMUX;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_AO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_AO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_BO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_BO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_CO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_CO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_DO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_DO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_AMUX;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_AO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_AO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_BMUX;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_BO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_BO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_CO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_DO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_DO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_AMUX;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_AO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_BMUX;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_BO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_CO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_CO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_DO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_DO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_AMUX;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_AO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_AO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_BMUX;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_BO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_CO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_CO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_DO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_AO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_AO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_BO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_BO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_CO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_DO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_DO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_AO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_BO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_BO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_CO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_CO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_DO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_DO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_AO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_AO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_BO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_BO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_CO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_CO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_DO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_DO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D_XOR;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A1;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A2;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A3;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A4;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_AMUX;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_AO5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_AO6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A_CY;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_A_XOR;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B1;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B2;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B3;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B4;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_BO5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_BO6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B_CY;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_B_XOR;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C1;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C2;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C3;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C4;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_CO5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_CO6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C_CY;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_C_XOR;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D1;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D2;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D3;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D4;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_DO5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_DO6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D_CY;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X20Y99_D_XOR;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A1;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A2;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A3;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A4;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_AO5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_AO6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A_CY;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_A_XOR;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B1;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B2;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B3;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B4;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_BO5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_BO6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B_CY;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_B_XOR;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C1;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C2;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C3;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C4;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_CO5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_CO6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C_CY;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_C_XOR;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D1;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D2;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D3;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D4;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_DO5;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_DO6;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D_CY;
  wire [0:0] CLBLM_R_X15Y99_SLICE_X21Y99_D_XOR;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A1;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A2;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A3;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A4;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_AO5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_AO6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A_CY;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_A_XOR;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B1;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B2;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B3;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B4;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_BO5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_BO6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B_CY;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_B_XOR;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C1;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C2;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C3;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C4;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_CO5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_CO6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C_CY;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_C_XOR;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D1;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D2;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D3;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D4;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_DO5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_DO6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D_CY;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X56Y111_D_XOR;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A1;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A2;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A3;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A4;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_AO5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_AO6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A_CY;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_A_XOR;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B1;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B2;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B3;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B4;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_BO5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_BO6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B_CY;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_B_XOR;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C1;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C2;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C3;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C4;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_CO5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_CO6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C_CY;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_C_XOR;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D1;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D2;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D3;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D4;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_DO5;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_DO6;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D_CY;
  wire [0:0] CLBLM_R_X37Y111_SLICE_X57Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_AO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_AO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_BO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_BO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_CO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_CO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_DO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_DO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_AO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_AO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_BO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_BO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_CO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_CO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_DO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_DO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_AO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_AO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_BO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_BO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_CO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_CO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_DO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_DO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_AO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_AO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_BO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_BO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_CO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_CO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_DO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_DO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_I;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_I;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y200_IOB_X0Y200_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_SING_X0Y99_IOB_X0Y99_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_I;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y81_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y82_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y83_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y84_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y85_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y86_I;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y87_I;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y88_I;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y89_I;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y90_I;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y91_I;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y92_I;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y93_I;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y94_I;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y95_I;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y96_I;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y97_I;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y98_I;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_D;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_O;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_D1;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_OQ;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_T1;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_SING_X0Y99_ILOGIC_X0Y99_D;
  wire [0:0] LIOI3_SING_X0Y99_ILOGIC_X0Y99_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_O;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y86_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y86_O;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y89_D;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y89_O;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y90_D;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y90_O;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y91_D;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y91_O;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y92_D;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y92_O;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y95_D;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y95_O;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y96_D;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y96_O;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y97_D;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y97_O;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y98_D;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y98_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_I;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_SING_X105Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_SING_X105Y99_IOB_X1Y99_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_I;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_I;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_I;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_I;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_I;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_I;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_I;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_I;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_I;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_I;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_I;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_I;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_I;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_I;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_I;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_I;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_I;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_I;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_I;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_I;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_I;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y53_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y54_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y56_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y57_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y59_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y60_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y62_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y63_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y64_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y65_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y66_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y67_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y68_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y69_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y70_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y71_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y72_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y73_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y74_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y77_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y78_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y79_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y80_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y81_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y82_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y83_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y84_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y85_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y86_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y87_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y88_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y89_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y90_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y91_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y92_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y93_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y94_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y95_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y96_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y97_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y98_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_SING_X105Y150_ILOGIC_X1Y150_D;
  wire [0:0] RIOI3_SING_X105Y150_ILOGIC_X1Y150_O;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y151_D;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y151_O;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y152_D;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y152_O;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y153_D;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y153_O;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y154_D;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y154_O;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y155_D;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y155_O;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y156_D;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y156_O;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y159_D;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y159_O;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y160_D;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y160_O;
  wire [0:0] RIOI3_X105Y161_ILOGIC_X1Y161_D;
  wire [0:0] RIOI3_X105Y161_ILOGIC_X1Y161_O;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y165_D;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y165_O;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y166_D;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y166_O;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y167_D;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y167_O;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y168_D;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y168_O;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y171_D;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y171_O;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y172_D;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y172_O;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_TQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_TQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y101_SLICE_X0Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y101_SLICE_X0Y101_DO5),
.O6(CLBLL_L_X2Y101_SLICE_X0Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005000400050004)
  ) CLBLL_L_X2Y101_SLICE_X0Y101_CLUT (
.I0(LIOB33_X0Y55_IOB_X0Y55_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y101_SLICE_X0Y101_CO5),
.O6(CLBLL_L_X2Y101_SLICE_X0Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffa)
  ) CLBLL_L_X2Y101_SLICE_X0Y101_BLUT (
.I0(LIOB33_X0Y59_IOB_X0Y60_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y78_I),
.I3(LIOB33_X0Y55_IOB_X0Y56_I),
.I4(CLBLL_L_X2Y101_SLICE_X0Y101_AO6),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLL_L_X2Y101_SLICE_X0Y101_BO5),
.O6(CLBLL_L_X2Y101_SLICE_X0Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffdffffffff)
  ) CLBLL_L_X2Y101_SLICE_X0Y101_ALUT (
.I0(LIOB33_X0Y63_IOB_X0Y63_I),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(LIOB33_X0Y75_IOB_X0Y75_I),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(LIOB33_X0Y71_IOB_X0Y72_I),
.I5(LIOB33_X0Y53_IOB_X0Y54_I),
.O5(CLBLL_L_X2Y101_SLICE_X0Y101_AO5),
.O6(CLBLL_L_X2Y101_SLICE_X0Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y101_SLICE_X1Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y101_SLICE_X1Y101_DO5),
.O6(CLBLL_L_X2Y101_SLICE_X1Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y101_SLICE_X1Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y101_SLICE_X1Y101_CO5),
.O6(CLBLL_L_X2Y101_SLICE_X1Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y101_SLICE_X1Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y101_SLICE_X1Y101_BO5),
.O6(CLBLL_L_X2Y101_SLICE_X1Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y101_SLICE_X1Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y101_SLICE_X1Y101_AO5),
.O6(CLBLL_L_X2Y101_SLICE_X1Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X0Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X0Y136_DO5),
.O6(CLBLL_L_X2Y136_SLICE_X0Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X0Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X0Y136_CO5),
.O6(CLBLL_L_X2Y136_SLICE_X0Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f00000)
  ) CLBLL_L_X2Y136_SLICE_X0Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(1'b1),
.I4(LIOB33_X0Y135_IOB_X0Y136_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X0Y136_BO5),
.O6(CLBLL_L_X2Y136_SLICE_X0Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLL_L_X2Y136_SLICE_X0Y136_ALUT (
.I0(LIOB33_X0Y137_IOB_X0Y138_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y67_IOB_X0Y67_I),
.I3(LIOB33_X0Y135_IOB_X0Y135_I),
.I4(LIOB33_X0Y135_IOB_X0Y136_I),
.I5(LIOB33_X0Y137_IOB_X0Y137_I),
.O5(CLBLL_L_X2Y136_SLICE_X0Y136_AO5),
.O6(CLBLL_L_X2Y136_SLICE_X0Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X1Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X1Y136_DO5),
.O6(CLBLL_L_X2Y136_SLICE_X1Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X1Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X1Y136_CO5),
.O6(CLBLL_L_X2Y136_SLICE_X1Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X1Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X1Y136_BO5),
.O6(CLBLL_L_X2Y136_SLICE_X1Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X1Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X1Y136_AO5),
.O6(CLBLL_L_X2Y136_SLICE_X1Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777ffffa0a0a0a0)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_ALUT (
.I0(LIOB33_X0Y75_IOB_X0Y76_I),
.I1(LIOB33_X0Y89_IOB_X0Y89_I),
.I2(LIOB33_X0Y145_IOB_X0Y146_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X0Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X0Y173_DO5),
.O6(CLBLL_L_X2Y173_SLICE_X0Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X0Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X0Y173_CO5),
.O6(CLBLL_L_X2Y173_SLICE_X0Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X0Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X0Y173_BO5),
.O6(CLBLL_L_X2Y173_SLICE_X0Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00a00000000000)
  ) CLBLL_L_X2Y173_SLICE_X0Y173_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y145_I),
.I1(1'b1),
.I2(LIOB33_X0Y173_IOB_X0Y173_I),
.I3(LIOB33_X0Y75_IOB_X0Y76_I),
.I4(LIOB33_X0Y171_IOB_X0Y172_I),
.I5(LIOB33_X0Y89_IOB_X0Y89_I),
.O5(CLBLL_L_X2Y173_SLICE_X0Y173_AO5),
.O6(CLBLL_L_X2Y173_SLICE_X0Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X1Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X1Y173_DO5),
.O6(CLBLL_L_X2Y173_SLICE_X1Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X1Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X1Y173_CO5),
.O6(CLBLL_L_X2Y173_SLICE_X1Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X1Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X1Y173_BO5),
.O6(CLBLL_L_X2Y173_SLICE_X1Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X1Y173_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X1Y173_AO5),
.O6(CLBLL_L_X2Y173_SLICE_X1Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y174_SLICE_X0Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y174_SLICE_X0Y174_DO5),
.O6(CLBLL_L_X2Y174_SLICE_X0Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y174_SLICE_X0Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y174_SLICE_X0Y174_CO5),
.O6(CLBLL_L_X2Y174_SLICE_X0Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00008800c0000000)
  ) CLBLL_L_X2Y174_SLICE_X0Y174_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_X0Y89_IOB_X0Y89_I),
.I2(LIOB33_X0Y171_IOB_X0Y171_I),
.I3(LIOB33_X0Y75_IOB_X0Y76_I),
.I4(LIOB33_X0Y145_IOB_X0Y145_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y174_SLICE_X0Y174_BO5),
.O6(CLBLL_L_X2Y174_SLICE_X0Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0000000f000f000)
  ) CLBLL_L_X2Y174_SLICE_X0Y174_ALUT (
.I0(LIOB33_X0Y173_IOB_X0Y174_I),
.I1(LIOB33_X0Y97_IOB_X0Y98_I),
.I2(LIOB33_X0Y89_IOB_X0Y89_I),
.I3(LIOB33_X0Y75_IOB_X0Y76_I),
.I4(LIOB33_X0Y145_IOB_X0Y145_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y174_SLICE_X0Y174_AO5),
.O6(CLBLL_L_X2Y174_SLICE_X0Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y174_SLICE_X1Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y174_SLICE_X1Y174_DO5),
.O6(CLBLL_L_X2Y174_SLICE_X1Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y174_SLICE_X1Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y174_SLICE_X1Y174_CO5),
.O6(CLBLL_L_X2Y174_SLICE_X1Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y174_SLICE_X1Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y174_SLICE_X1Y174_BO5),
.O6(CLBLL_L_X2Y174_SLICE_X1Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y174_SLICE_X1Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y174_SLICE_X1Y174_AO5),
.O6(CLBLL_L_X2Y174_SLICE_X1Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X0Y175_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X0Y175_DO5),
.O6(CLBLL_L_X2Y175_SLICE_X0Y175_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X0Y175_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X0Y175_CO5),
.O6(CLBLL_L_X2Y175_SLICE_X0Y175_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X0Y175_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X0Y175_BO5),
.O6(CLBLL_L_X2Y175_SLICE_X0Y175_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f00000)
  ) CLBLL_L_X2Y175_SLICE_X0Y175_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y137_IOB_X0Y138_I),
.I3(1'b1),
.I4(LIOB33_X0Y135_IOB_X0Y135_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X0Y175_AO5),
.O6(CLBLL_L_X2Y175_SLICE_X0Y175_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X1Y175_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X1Y175_DO5),
.O6(CLBLL_L_X2Y175_SLICE_X1Y175_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X1Y175_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X1Y175_CO5),
.O6(CLBLL_L_X2Y175_SLICE_X1Y175_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X1Y175_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X1Y175_BO5),
.O6(CLBLL_L_X2Y175_SLICE_X1Y175_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X1Y175_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X1Y175_AO5),
.O6(CLBLL_L_X2Y175_SLICE_X1Y175_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X160Y125_DO5),
.O6(CLBLL_L_X102Y125_SLICE_X160Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X160Y125_CO5),
.O6(CLBLL_L_X102Y125_SLICE_X160Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X160Y125_BO5),
.O6(CLBLL_L_X102Y125_SLICE_X160Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X160Y125_AO5),
.O6(CLBLL_L_X102Y125_SLICE_X160Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X161Y125_DO5),
.O6(CLBLL_L_X102Y125_SLICE_X161Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X161Y125_CO5),
.O6(CLBLL_L_X102Y125_SLICE_X161Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc00fc00cc00dc00)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I1(CLBLM_R_X103Y125_SLICE_X163Y125_AO6),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I3(CLBLL_R_X81Y124_SLICE_X126Y124_AO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I5(CLBLM_R_X15Y114_SLICE_X20Y114_AO5),
.O5(CLBLL_L_X102Y125_SLICE_X161Y125_BO5),
.O6(CLBLL_L_X102Y125_SLICE_X161Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0000ccdc0000)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_ALUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I1(CLBLM_R_X103Y125_SLICE_X163Y125_AO6),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I4(CLBLL_R_X81Y122_SLICE_X126Y122_CO6),
.I5(CLBLM_R_X15Y114_SLICE_X20Y114_AO5),
.O5(CLBLL_L_X102Y125_SLICE_X161Y125_AO5),
.O6(CLBLL_L_X102Y125_SLICE_X161Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y111_SLICE_X126Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y111_SLICE_X126Y111_DO5),
.O6(CLBLL_R_X81Y111_SLICE_X126Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y111_SLICE_X126Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y111_SLICE_X126Y111_CO5),
.O6(CLBLL_R_X81Y111_SLICE_X126Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300003331)
  ) CLBLL_R_X81Y111_SLICE_X126Y111_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I1(LIOB33_X0Y157_IOB_X0Y157_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(LIOB33_X0Y165_IOB_X0Y165_I),
.I4(LIOB33_X0Y157_IOB_X0Y158_I),
.I5(CLBLM_R_X13Y112_SLICE_X19Y112_DO6),
.O5(CLBLL_R_X81Y111_SLICE_X126Y111_BO5),
.O6(CLBLL_R_X81Y111_SLICE_X126Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ff000000fd)
  ) CLBLL_R_X81Y111_SLICE_X126Y111_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I1(LIOB33_X0Y165_IOB_X0Y165_I),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(LIOB33_X0Y153_IOB_X0Y154_I),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(CLBLM_R_X13Y112_SLICE_X19Y112_DO6),
.O5(CLBLL_R_X81Y111_SLICE_X126Y111_AO5),
.O6(CLBLL_R_X81Y111_SLICE_X126Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y111_SLICE_X127Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y111_SLICE_X127Y111_DO5),
.O6(CLBLL_R_X81Y111_SLICE_X127Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y111_SLICE_X127Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y111_SLICE_X127Y111_CO5),
.O6(CLBLL_R_X81Y111_SLICE_X127Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y111_SLICE_X127Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y111_SLICE_X127Y111_BO5),
.O6(CLBLL_R_X81Y111_SLICE_X127Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y111_SLICE_X127Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y111_SLICE_X127Y111_AO5),
.O6(CLBLL_R_X81Y111_SLICE_X127Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y122_SLICE_X126Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y122_SLICE_X126Y122_DO5),
.O6(CLBLL_R_X81Y122_SLICE_X126Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ff000000ff)
  ) CLBLL_R_X81Y122_SLICE_X126Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y157_IOB_X0Y157_I),
.I4(LIOB33_X0Y157_IOB_X0Y158_I),
.I5(1'b1),
.O5(CLBLL_R_X81Y122_SLICE_X126Y122_CO5),
.O6(CLBLL_R_X81Y122_SLICE_X126Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055555554)
  ) CLBLL_R_X81Y122_SLICE_X126Y122_BLUT (
.I0(LIOB33_X0Y157_IOB_X0Y158_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(LIOB33_X0Y155_IOB_X0Y155_I),
.I3(RIOB33_X105Y155_IOB_X1Y155_I),
.I4(CLBLM_R_X13Y110_SLICE_X19Y110_CO6),
.I5(LIOB33_X0Y157_IOB_X0Y157_I),
.O5(CLBLL_R_X81Y122_SLICE_X126Y122_BO5),
.O6(CLBLL_R_X81Y122_SLICE_X126Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505050504)
  ) CLBLL_R_X81Y122_SLICE_X126Y122_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(RIOB33_X105Y155_IOB_X1Y155_I),
.I4(LIOB33_X0Y155_IOB_X0Y155_I),
.I5(CLBLM_R_X13Y110_SLICE_X19Y110_CO6),
.O5(CLBLL_R_X81Y122_SLICE_X126Y122_AO5),
.O6(CLBLL_R_X81Y122_SLICE_X126Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y122_SLICE_X127Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y122_SLICE_X127Y122_DO5),
.O6(CLBLL_R_X81Y122_SLICE_X127Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y122_SLICE_X127Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y122_SLICE_X127Y122_CO5),
.O6(CLBLL_R_X81Y122_SLICE_X127Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y122_SLICE_X127Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y122_SLICE_X127Y122_BO5),
.O6(CLBLL_R_X81Y122_SLICE_X127Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y122_SLICE_X127Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y122_SLICE_X127Y122_AO5),
.O6(CLBLL_R_X81Y122_SLICE_X127Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y124_SLICE_X126Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y124_SLICE_X126Y124_DO5),
.O6(CLBLL_R_X81Y124_SLICE_X126Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y124_SLICE_X126Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y124_SLICE_X126Y124_CO5),
.O6(CLBLL_R_X81Y124_SLICE_X126Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y124_SLICE_X126Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y124_SLICE_X126Y124_BO5),
.O6(CLBLL_R_X81Y124_SLICE_X126Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505050505)
  ) CLBLL_R_X81Y124_SLICE_X126Y124_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(1'b1),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y124_SLICE_X126Y124_AO5),
.O6(CLBLL_R_X81Y124_SLICE_X126Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y124_SLICE_X127Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y124_SLICE_X127Y124_DO5),
.O6(CLBLL_R_X81Y124_SLICE_X127Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y124_SLICE_X127Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y124_SLICE_X127Y124_CO5),
.O6(CLBLL_R_X81Y124_SLICE_X127Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y124_SLICE_X127Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y124_SLICE_X127Y124_BO5),
.O6(CLBLL_R_X81Y124_SLICE_X127Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X81Y124_SLICE_X127Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X81Y124_SLICE_X127Y124_AO5),
.O6(CLBLL_R_X81Y124_SLICE_X127Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddffdfff99ff9aff)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y95_IOB_X0Y96_I),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.I4(LIOB33_X0Y77_IOB_X0Y78_I),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f000003)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeccffcffe)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y75_IOB_X0Y75_I),
.I5(LIOB33_X0Y95_IOB_X0Y96_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fa00faccfeccfe)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y75_IOB_X0Y75_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff5f00ff00f0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(1'b1),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y77_IOB_X0Y78_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff3b00000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y78_I),
.I3(RIOB33_X105Y167_IOB_X1Y168_I),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffbf0f0f)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(LIOB33_X0Y75_IOB_X0Y75_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I5(RIOB33_X105Y169_IOB_X1Y169_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000004)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0f0fefff)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0f0f000f0b0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff20ff2)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaaeaaafaaaeaa)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(RIOB33_X105Y165_IOB_X1Y166_I),
.I1(LIOB33_X0Y151_IOB_X0Y151_I),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f5f700000000)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I2(LIOB33_X0Y129_IOB_X0Y130_I),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005555f3f0f2f0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(LIOB33_X0Y129_IOB_X0Y130_I),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(LIOB33_X0Y151_IOB_X0Y151_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y93_IOB_X0Y93_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fffffffffffe)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_ALUT (
.I0(LIOB33_X0Y87_IOB_X0Y88_I),
.I1(LIOB33_X0Y91_IOB_X0Y91_I),
.I2(LIOB33_X0Y85_IOB_X0Y86_I),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X30Y111_SLICE_X44Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X30Y111_SLICE_X44Y111_DO5),
.O6(CLBLM_L_X30Y111_SLICE_X44Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X30Y111_SLICE_X44Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X30Y111_SLICE_X44Y111_CO5),
.O6(CLBLM_L_X30Y111_SLICE_X44Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000fffe)
  ) CLBLM_L_X30Y111_SLICE_X44Y111_BLUT (
.I0(CLBLM_R_X13Y113_SLICE_X19Y113_CO6),
.I1(LIOB33_X0Y163_IOB_X0Y163_I),
.I2(LIOB33_X0Y163_IOB_X0Y164_I),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(LIOB33_X0Y157_IOB_X0Y158_I),
.O5(CLBLM_L_X30Y111_SLICE_X44Y111_BO5),
.O6(CLBLM_L_X30Y111_SLICE_X44Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000fffe)
  ) CLBLM_L_X30Y111_SLICE_X44Y111_ALUT (
.I0(LIOB33_X0Y163_IOB_X0Y164_I),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_CO6),
.I2(LIOB33_X0Y163_IOB_X0Y163_I),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(LIOB33_X0Y153_IOB_X0Y154_I),
.O5(CLBLM_L_X30Y111_SLICE_X44Y111_AO5),
.O6(CLBLM_L_X30Y111_SLICE_X44Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X30Y111_SLICE_X45Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X30Y111_SLICE_X45Y111_DO5),
.O6(CLBLM_L_X30Y111_SLICE_X45Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X30Y111_SLICE_X45Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X30Y111_SLICE_X45Y111_CO5),
.O6(CLBLM_L_X30Y111_SLICE_X45Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X30Y111_SLICE_X45Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X30Y111_SLICE_X45Y111_BO5),
.O6(CLBLM_L_X30Y111_SLICE_X45Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X30Y111_SLICE_X45Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X30Y111_SLICE_X45Y111_AO5),
.O6(CLBLM_L_X30Y111_SLICE_X45Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y121_SLICE_X70Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y121_SLICE_X70Y121_DO5),
.O6(CLBLM_L_X46Y121_SLICE_X70Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y121_SLICE_X70Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y121_SLICE_X70Y121_CO5),
.O6(CLBLM_L_X46Y121_SLICE_X70Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaafaffffeefe)
  ) CLBLM_L_X46Y121_SLICE_X70Y121_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X15Y110_SLICE_X20Y110_BO6),
.I2(LIOB33_X0Y175_IOB_X0Y176_I),
.I3(LIOB33_X0Y159_IOB_X0Y160_I),
.I4(RIOB33_X105Y119_IOB_X1Y120_I),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_CO6),
.O5(CLBLM_L_X46Y121_SLICE_X70Y121_BO5),
.O6(CLBLM_L_X46Y121_SLICE_X70Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaafaffffeefe)
  ) CLBLM_L_X46Y121_SLICE_X70Y121_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X15Y110_SLICE_X20Y110_BO6),
.I2(LIOB33_X0Y175_IOB_X0Y176_I),
.I3(LIOB33_X0Y159_IOB_X0Y160_I),
.I4(LIOB33_X0Y161_IOB_X0Y162_I),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_CO6),
.O5(CLBLM_L_X46Y121_SLICE_X70Y121_AO5),
.O6(CLBLM_L_X46Y121_SLICE_X70Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y121_SLICE_X71Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y121_SLICE_X71Y121_DO5),
.O6(CLBLM_L_X46Y121_SLICE_X71Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y121_SLICE_X71Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y121_SLICE_X71Y121_CO5),
.O6(CLBLM_L_X46Y121_SLICE_X71Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y121_SLICE_X71Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y121_SLICE_X71Y121_BO5),
.O6(CLBLM_L_X46Y121_SLICE_X71Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y121_SLICE_X71Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y121_SLICE_X71Y121_AO5),
.O6(CLBLM_L_X46Y121_SLICE_X71Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y142_SLICE_X70Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y142_SLICE_X70Y142_DO5),
.O6(CLBLM_L_X46Y142_SLICE_X70Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y142_SLICE_X70Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y142_SLICE_X70Y142_CO5),
.O6(CLBLM_L_X46Y142_SLICE_X70Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y142_SLICE_X70Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y142_SLICE_X70Y142_BO5),
.O6(CLBLM_L_X46Y142_SLICE_X70Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0ffff)
  ) CLBLM_L_X46Y142_SLICE_X70Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y159_IOB_X0Y160_I),
.I3(1'b1),
.I4(LIOB33_X0Y177_IOB_X0Y177_I),
.I5(1'b1),
.O5(CLBLM_L_X46Y142_SLICE_X70Y142_AO5),
.O6(CLBLM_L_X46Y142_SLICE_X70Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y142_SLICE_X71Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y142_SLICE_X71Y142_DO5),
.O6(CLBLM_L_X46Y142_SLICE_X71Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y142_SLICE_X71Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y142_SLICE_X71Y142_CO5),
.O6(CLBLM_L_X46Y142_SLICE_X71Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y142_SLICE_X71Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y142_SLICE_X71Y142_BO5),
.O6(CLBLM_L_X46Y142_SLICE_X71Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y142_SLICE_X71Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y142_SLICE_X71Y142_AO5),
.O6(CLBLM_L_X46Y142_SLICE_X71Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y119_SLICE_X76Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y119_SLICE_X76Y119_DO5),
.O6(CLBLM_L_X50Y119_SLICE_X76Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y119_SLICE_X76Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y119_SLICE_X76Y119_CO5),
.O6(CLBLM_L_X50Y119_SLICE_X76Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y119_SLICE_X76Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y119_SLICE_X76Y119_BO5),
.O6(CLBLM_L_X50Y119_SLICE_X76Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfcfffafffa)
  ) CLBLM_L_X50Y119_SLICE_X76Y119_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(LIOB33_X0Y175_IOB_X0Y175_I),
.I2(CLBLM_R_X15Y113_SLICE_X21Y113_DO6),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_L_X50Y119_SLICE_X76Y119_AO5),
.O6(CLBLM_L_X50Y119_SLICE_X76Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y119_SLICE_X77Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y119_SLICE_X77Y119_DO5),
.O6(CLBLM_L_X50Y119_SLICE_X77Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y119_SLICE_X77Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y119_SLICE_X77Y119_CO5),
.O6(CLBLM_L_X50Y119_SLICE_X77Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y119_SLICE_X77Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y119_SLICE_X77Y119_BO5),
.O6(CLBLM_L_X50Y119_SLICE_X77Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X50Y119_SLICE_X77Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X50Y119_SLICE_X77Y119_AO5),
.O6(CLBLM_L_X50Y119_SLICE_X77Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X120Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X120Y119_DO5),
.O6(CLBLM_L_X78Y119_SLICE_X120Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X120Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X120Y119_CO5),
.O6(CLBLM_L_X78Y119_SLICE_X120Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X120Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X120Y119_BO5),
.O6(CLBLM_L_X78Y119_SLICE_X120Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X120Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X120Y119_AO5),
.O6(CLBLM_L_X78Y119_SLICE_X120Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5d0000ff000000)
  ) CLBLM_L_X78Y119_SLICE_X121Y119_DLUT (
.I0(CLBLM_R_X15Y114_SLICE_X20Y114_BO5),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I3(CLBLM_L_X50Y119_SLICE_X76Y119_AO5),
.I4(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O5(CLBLM_L_X78Y119_SLICE_X121Y119_DO5),
.O6(CLBLM_L_X78Y119_SLICE_X121Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc4ccc44cc00cc00)
  ) CLBLM_L_X78Y119_SLICE_X121Y119_CLUT (
.I0(CLBLM_R_X15Y114_SLICE_X20Y114_BO5),
.I1(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I3(CLBLM_L_X50Y119_SLICE_X76Y119_AO5),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O5(CLBLM_L_X78Y119_SLICE_X121Y119_CO5),
.O6(CLBLM_L_X78Y119_SLICE_X121Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a8a8a8a0a0a8a8)
  ) CLBLM_L_X78Y119_SLICE_X121Y119_BLUT (
.I0(CLBLL_R_X81Y122_SLICE_X126Y122_CO6),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(CLBLM_L_X50Y119_SLICE_X76Y119_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I4(CLBLM_R_X15Y114_SLICE_X20Y114_BO5),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.O5(CLBLM_L_X78Y119_SLICE_X121Y119_BO5),
.O6(CLBLM_L_X78Y119_SLICE_X121Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f020a0f0f000a0)
  ) CLBLM_L_X78Y119_SLICE_X121Y119_ALUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I2(CLBLL_R_X81Y124_SLICE_X126Y124_AO6),
.I3(CLBLM_R_X15Y114_SLICE_X20Y114_BO5),
.I4(CLBLM_L_X50Y119_SLICE_X76Y119_AO6),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.O5(CLBLM_L_X78Y119_SLICE_X121Y119_AO5),
.O6(CLBLM_L_X78Y119_SLICE_X121Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y125_SLICE_X120Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y125_SLICE_X120Y125_DO5),
.O6(CLBLM_L_X78Y125_SLICE_X120Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y125_SLICE_X120Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y125_SLICE_X120Y125_CO5),
.O6(CLBLM_L_X78Y125_SLICE_X120Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y125_SLICE_X120Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y125_SLICE_X120Y125_BO5),
.O6(CLBLM_L_X78Y125_SLICE_X120Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y125_SLICE_X120Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y125_SLICE_X120Y125_AO5),
.O6(CLBLM_L_X78Y125_SLICE_X120Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f5007500)
  ) CLBLM_L_X78Y125_SLICE_X121Y125_DLUT (
.I0(CLBLM_L_X46Y142_SLICE_X70Y142_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I3(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I5(CLBLM_L_X46Y121_SLICE_X70Y121_BO6),
.O5(CLBLM_L_X78Y125_SLICE_X121Y125_DO5),
.O6(CLBLM_L_X78Y125_SLICE_X121Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccc4c444c4)
  ) CLBLM_L_X78Y125_SLICE_X121Y125_CLUT (
.I0(CLBLM_L_X46Y142_SLICE_X70Y142_AO6),
.I1(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I5(CLBLM_L_X46Y121_SLICE_X70Y121_BO6),
.O5(CLBLM_L_X78Y125_SLICE_X121Y125_CO5),
.O6(CLBLM_L_X78Y125_SLICE_X121Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf080f0f0f0c0f0f0)
  ) CLBLM_L_X78Y125_SLICE_X121Y125_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(CLBLL_R_X81Y122_SLICE_X126Y122_CO6),
.I3(CLBLM_L_X46Y121_SLICE_X70Y121_AO6),
.I4(CLBLM_L_X46Y142_SLICE_X70Y142_AO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.O5(CLBLM_L_X78Y125_SLICE_X121Y125_BO5),
.O6(CLBLM_L_X78Y125_SLICE_X121Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008f00ff00cf00)
  ) CLBLM_L_X78Y125_SLICE_X121Y125_ALUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(CLBLM_L_X46Y142_SLICE_X70Y142_AO6),
.I3(CLBLL_R_X81Y124_SLICE_X126Y124_AO6),
.I4(CLBLM_L_X46Y121_SLICE_X70Y121_AO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.O5(CLBLM_L_X78Y125_SLICE_X121Y125_AO5),
.O6(CLBLM_L_X78Y125_SLICE_X121Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X144Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X144Y125_DO5),
.O6(CLBLM_L_X92Y125_SLICE_X144Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X144Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X144Y125_CO5),
.O6(CLBLM_L_X92Y125_SLICE_X144Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300000003030000)
  ) CLBLM_L_X92Y125_SLICE_X144Y125_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y141_IOB_X0Y142_I),
.I2(LIOB33_X0Y143_IOB_X0Y143_I),
.I3(CLBLM_R_X103Y122_SLICE_X163Y122_AO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.O6(CLBLM_L_X92Y125_SLICE_X144Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300000003030000)
  ) CLBLM_L_X92Y125_SLICE_X144Y125_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y139_IOB_X0Y140_I),
.I2(LIOB33_X0Y141_IOB_X0Y141_I),
.I3(CLBLM_R_X103Y122_SLICE_X163Y122_AO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.O6(CLBLM_L_X92Y125_SLICE_X144Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X145Y125_DO5),
.O6(CLBLM_L_X92Y125_SLICE_X145Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X145Y125_CO5),
.O6(CLBLM_L_X92Y125_SLICE_X145Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X145Y125_BO5),
.O6(CLBLM_L_X92Y125_SLICE_X145Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X145Y125_AO5),
.O6(CLBLM_L_X92Y125_SLICE_X145Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X148Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X148Y122_DO5),
.O6(CLBLM_L_X94Y122_SLICE_X148Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X148Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X148Y122_CO5),
.O6(CLBLM_L_X94Y122_SLICE_X148Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa88aa8aaa00aa00)
  ) CLBLM_L_X94Y122_SLICE_X148Y122_BLUT (
.I0(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I3(CLBLM_R_X93Y116_SLICE_X147Y116_AO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O5(CLBLM_L_X94Y122_SLICE_X148Y122_BO5),
.O6(CLBLM_L_X94Y122_SLICE_X148Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa88008a00)
  ) CLBLM_L_X94Y122_SLICE_X148Y122_ALUT (
.I0(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I3(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I5(CLBLM_R_X93Y116_SLICE_X147Y116_AO6),
.O5(CLBLM_L_X94Y122_SLICE_X148Y122_AO5),
.O6(CLBLM_L_X94Y122_SLICE_X148Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X149Y122_DO5),
.O6(CLBLM_L_X94Y122_SLICE_X149Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X149Y122_CO5),
.O6(CLBLM_L_X94Y122_SLICE_X149Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X149Y122_BO5),
.O6(CLBLM_L_X94Y122_SLICE_X149Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X149Y122_AO5),
.O6(CLBLM_L_X94Y122_SLICE_X149Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333300000004)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(CLBLM_R_X13Y109_SLICE_X18Y109_AO6),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I2(CLBLL_L_X2Y136_SLICE_X0Y136_AO6),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.I4(CLBLL_L_X2Y101_SLICE_X0Y101_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffff00)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y59_IOB_X0Y60_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(LIOB33_X0Y95_IOB_X0Y96_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff33337777)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y79_IOB_X0Y80_I),
.I5(LIOB33_X0Y95_IOB_X0Y96_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(CLBLL_L_X2Y101_SLICE_X0Y101_CO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h323232320000cdcd)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(LIOB33_X0Y57_IOB_X0Y57_I),
.I1(LIOB33_X0Y95_IOB_X0Y96_I),
.I2(LIOB33_X0Y55_IOB_X0Y56_I),
.I3(1'b1),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffddffddff)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y55_IOB_X0Y56_I),
.I2(1'b1),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(1'b1),
.I5(LIOB33_X0Y57_IOB_X0Y58_I),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000c00)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y79_IOB_X0Y80_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y75_IOB_X0Y75_I),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00dc00ff00ff00)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(RIOB33_X105Y161_IOB_X1Y161_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf30ff35bcfcccfcd)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa4410aaaa4410)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff3fffffff2)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y95_IOB_X0Y96_I),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he5e5e5eeafafafaa)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y77_IOB_X0Y78_I),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafafb0f0c0f0c)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y59_IOB_X0Y59_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020002000200030)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(LIOB33_X0Y95_IOB_X0Y96_I),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.I4(LIOB33_X0Y79_IOB_X0Y80_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf3fdf3fdf3fdfdf)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y79_IOB_X0Y80_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccc080000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffceeeefffe)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y79_IOB_X0Y80_I),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefefeffffffff)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f7ffffffffffff)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.I1(LIOB33_X0Y59_IOB_X0Y59_I),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I5(LIOB33_X0Y121_IOB_X0Y122_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33223322cccccfcf)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(LIOB33_X0Y65_IOB_X0Y65_I),
.I1(LIOB33_X0Y95_IOB_X0Y96_I),
.I2(LIOB33_X0Y73_IOB_X0Y74_I),
.I3(LIOB33_X0Y63_IOB_X0Y63_I),
.I4(LIOB33_X0Y71_IOB_X0Y72_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000003ff00ff00)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeeeaaaaaeeee)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f0000fe0f0000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaafaeeffeefe)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.I2(LIOB33_X0Y71_IOB_X0Y72_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y73_IOB_X0Y74_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040004000)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff6fffffffff)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I5(LIOB33_X0Y139_IOB_X0Y139_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f01010000e0e0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(LIOB33_X0Y59_IOB_X0Y60_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(1'b1),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550011ffff5577)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(LIOB33_X0Y63_IOB_X0Y63_I),
.I2(1'b1),
.I3(LIOB33_X0Y65_IOB_X0Y65_I),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000a000a00)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(1'b1),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(1'b1),
.I5(LIOB33_X0Y71_IOB_X0Y72_I),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffffaa88)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y151_IOB_X0Y151_I),
.I2(1'b1),
.I3(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I4(RIOB33_X105Y169_IOB_X1Y170_I),
.I5(LIOB33_X0Y71_IOB_X0Y72_I),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c0c400000000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y59_IOB_X0Y60_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffff0000c0c4)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(LIOB33_X0Y59_IOB_X0Y59_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffff7ff)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(LIOB33_X0Y119_IOB_X0Y119_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I5(LIOB33_X0Y59_IOB_X0Y60_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y78_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f30f0ca0a2)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(LIOB33_X0Y55_IOB_X0Y55_I),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(LIOB33_X0Y119_IOB_X0Y119_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff88ff88ff)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(LIOB33_X0Y119_IOB_X0Y119_I),
.I1(LIOB33_X0Y53_IOB_X0Y54_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(LIOB33_X0Y59_IOB_X0Y60_I),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff80ff82ff80ff82)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y78_I),
.I3(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333303033333030)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y95_IOB_X0Y95_I),
.I2(LIOB33_X0Y85_IOB_X0Y86_I),
.I3(1'b1),
.I4(LIOB33_X0Y87_IOB_X0Y87_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_DO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcfdffff)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X13Y110_SLICE_X19Y110_AO5),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_CO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff33333332)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_BLUT (
.I0(LIOB33_X0Y87_IOB_X0Y87_I),
.I1(LIOB33_X0Y95_IOB_X0Y95_I),
.I2(LIOB33_X0Y91_IOB_X0Y91_I),
.I3(LIOB33_X0Y85_IOB_X0Y86_I),
.I4(LIOB33_X0Y91_IOB_X0Y92_I),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_AO6),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_BO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff3fff2)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_ALUT (
.I0(LIOB33_X0Y87_IOB_X0Y88_I),
.I1(LIOB33_X0Y95_IOB_X0Y95_I),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_R_X13Y109_SLICE_X18Y109_BO6),
.I4(LIOB33_X0Y89_IOB_X0Y90_I),
.I5(CLBLM_R_X13Y109_SLICE_X18Y109_CO6),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_AO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_DO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_CO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_BO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_AO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_DO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_CO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_BO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_AO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_DO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4c4c4ccc0c0c0cc)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_CLUT (
.I0(LIOB33_X0Y131_IOB_X0Y132_I),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I5(CLBLM_R_X13Y110_SLICE_X19Y110_BO6),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_CO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccff32323232)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_BLUT (
.I0(LIOB33_X0Y93_IOB_X0Y94_I),
.I1(LIOB33_X0Y95_IOB_X0Y95_I),
.I2(LIOB33_X0Y93_IOB_X0Y93_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333303030303)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_AO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_DO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_CO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0f0f0f0e)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_BLUT (
.I0(LIOB33_X0Y91_IOB_X0Y91_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(LIOB33_X0Y91_IOB_X0Y92_I),
.I5(LIOB33_X0Y125_IOB_X0Y125_I),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_ALUT (
.I0(CLBLM_R_X13Y112_SLICE_X18Y112_AO5),
.I1(CLBLM_R_X13Y110_SLICE_X19Y110_BO6),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_BO6),
.I4(LIOB33_X0Y131_IOB_X0Y132_I),
.I5(LIOB33_X0Y131_IOB_X0Y131_I),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_AO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_DO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_CO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_BO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fc00fc00ff00aa)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_ALUT (
.I0(LIOB33_X0Y91_IOB_X0Y91_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y95_IOB_X0Y95_I),
.I4(LIOB33_X0Y91_IOB_X0Y92_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_AO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ffabffabff)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_DLUT (
.I0(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I1(LIOB33_X0Y131_IOB_X0Y132_I),
.I2(CLBLM_R_X13Y110_SLICE_X19Y110_BO6),
.I3(CLBLM_R_X13Y112_SLICE_X18Y112_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y131_IOB_X0Y131_I),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_DO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbfffff)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_CLUT (
.I0(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(LIOB33_X0Y129_IOB_X0Y129_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_X0Y131_IOB_X0Y131_I),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_BO6),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_CO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefcdeecceecceecc)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y93_IOB_X0Y93_I),
.I3(LIOB33_X0Y69_IOB_X0Y70_I),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_BO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33303330bbbabbba)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_ALUT (
.I0(LIOB33_X0Y129_IOB_X0Y129_I),
.I1(LIOB33_X0Y95_IOB_X0Y95_I),
.I2(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_AO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8c8c8c8c8c8ccc8c)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_DLUT (
.I0(RIOB33_X105Y163_IOB_X1Y163_I),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(CLBLM_R_X13Y112_SLICE_X18Y112_DO6),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_DO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f1f10f0f0f0e)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y131_IOB_X0Y131_I),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_CO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffffffffffff)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_BLUT (
.I0(LIOB33_X0Y129_IOB_X0Y129_I),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(LIOB33_X0Y93_IOB_X0Y93_I),
.I3(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(LIOB33_X0Y151_IOB_X0Y151_I),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_BO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I1(LIOB33_X0Y131_IOB_X0Y131_I),
.I2(CLBLM_R_X15Y111_SLICE_X21Y111_AO5),
.I3(CLBLM_R_X13Y112_SLICE_X19Y112_BO6),
.I4(CLBLM_R_X15Y110_SLICE_X20Y110_BO6),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_AO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_DO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_CO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_BO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0c000c00)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y131_IOB_X0Y131_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(1'b1),
.I5(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_AO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5e5f5a5affffffff)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_DLUT (
.I0(CLBLM_R_X13Y112_SLICE_X18Y112_AO6),
.I1(CLBLM_R_X13Y110_SLICE_X19Y110_BO6),
.I2(LIOB33_X0Y129_IOB_X0Y129_I),
.I3(CLBLM_R_X13Y113_SLICE_X19Y113_AO5),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_CO6),
.I5(CLBLM_R_X13Y113_SLICE_X19Y113_BO6),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_DO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5f400000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_CLUT (
.I0(CLBLM_R_X13Y113_SLICE_X19Y113_AO6),
.I1(CLBLM_R_X13Y110_SLICE_X19Y110_BO6),
.I2(RIOB33_X105Y171_IOB_X1Y171_I),
.I3(LIOB33_X0Y131_IOB_X0Y132_I),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_AO6),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_CO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcff3e3f3e3)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_BLUT (
.I0(LIOB33_X0Y129_IOB_X0Y129_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(LIOB33_X0Y131_IOB_X0Y131_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050505540404044)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_ALUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(LIOB33_X0Y131_IOB_X0Y132_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_AO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y99_SLICE_X20Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y99_SLICE_X20Y99_DO5),
.O6(CLBLM_R_X15Y99_SLICE_X20Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y99_SLICE_X20Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y99_SLICE_X20Y99_CO5),
.O6(CLBLM_R_X15Y99_SLICE_X20Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y99_SLICE_X20Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y99_SLICE_X20Y99_BO5),
.O6(CLBLM_R_X15Y99_SLICE_X20Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55505550aaafaaaf)
  ) CLBLM_R_X15Y99_SLICE_X20Y99_ALUT (
.I0(LIOB33_X0Y95_IOB_X0Y95_I),
.I1(1'b1),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y99_SLICE_X20Y99_AO5),
.O6(CLBLM_R_X15Y99_SLICE_X20Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y99_SLICE_X21Y99_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y99_SLICE_X21Y99_DO5),
.O6(CLBLM_R_X15Y99_SLICE_X21Y99_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y99_SLICE_X21Y99_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y99_SLICE_X21Y99_CO5),
.O6(CLBLM_R_X15Y99_SLICE_X21Y99_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y99_SLICE_X21Y99_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y99_SLICE_X21Y99_BO5),
.O6(CLBLM_R_X15Y99_SLICE_X21Y99_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y99_SLICE_X21Y99_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y99_SLICE_X21Y99_AO5),
.O6(CLBLM_R_X15Y99_SLICE_X21Y99_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y101_SLICE_X20Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X20Y101_DO5),
.O6(CLBLM_R_X15Y101_SLICE_X20Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y101_SLICE_X20Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X20Y101_CO5),
.O6(CLBLM_R_X15Y101_SLICE_X20Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y101_SLICE_X20Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X20Y101_BO5),
.O6(CLBLM_R_X15Y101_SLICE_X20Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55af507788738c)
  ) CLBLM_R_X15Y101_SLICE_X20Y101_ALUT (
.I0(LIOB33_X0Y95_IOB_X0Y95_I),
.I1(CLBLM_R_X15Y109_SLICE_X20Y109_AO5),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y85_IOB_X0Y85_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X20Y101_AO5),
.O6(CLBLM_R_X15Y101_SLICE_X20Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y101_SLICE_X21Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X21Y101_DO5),
.O6(CLBLM_R_X15Y101_SLICE_X21Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y101_SLICE_X21Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X21Y101_CO5),
.O6(CLBLM_R_X15Y101_SLICE_X21Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y101_SLICE_X21Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X21Y101_BO5),
.O6(CLBLM_R_X15Y101_SLICE_X21Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y101_SLICE_X21Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X21Y101_AO5),
.O6(CLBLM_R_X15Y101_SLICE_X21Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y109_SLICE_X20Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X20Y109_DO5),
.O6(CLBLM_R_X15Y109_SLICE_X20Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y109_SLICE_X20Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X20Y109_CO5),
.O6(CLBLM_R_X15Y109_SLICE_X20Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200660020006500)
  ) CLBLM_R_X15Y109_SLICE_X20Y109_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_X0Y95_IOB_X0Y95_I),
.I2(LIOB33_X0Y93_IOB_X0Y93_I),
.I3(CLBLM_R_X15Y99_SLICE_X20Y99_AO5),
.I4(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.I5(LIOB33_X0Y93_IOB_X0Y94_I),
.O5(CLBLM_R_X15Y109_SLICE_X20Y109_BO5),
.O6(CLBLM_R_X15Y109_SLICE_X20Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f2f2f3b9b9b9fc)
  ) CLBLM_R_X15Y109_SLICE_X20Y109_ALUT (
.I0(LIOB33_X0Y95_IOB_X0Y95_I),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.I3(LIOB33_X0Y93_IOB_X0Y93_I),
.I4(LIOB33_X0Y93_IOB_X0Y94_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X20Y109_AO5),
.O6(CLBLM_R_X15Y109_SLICE_X20Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y109_SLICE_X21Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X21Y109_DO5),
.O6(CLBLM_R_X15Y109_SLICE_X21Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y109_SLICE_X21Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X21Y109_CO5),
.O6(CLBLM_R_X15Y109_SLICE_X21Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y109_SLICE_X21Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X21Y109_BO5),
.O6(CLBLM_R_X15Y109_SLICE_X21Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y109_SLICE_X21Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X21Y109_AO5),
.O6(CLBLM_R_X15Y109_SLICE_X21Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800880000000000)
  ) CLBLM_R_X15Y110_SLICE_X20Y110_DLUT (
.I0(LIOB33_X0Y153_IOB_X0Y153_I),
.I1(LIOB33_X0Y161_IOB_X0Y161_I),
.I2(CLBLM_R_X15Y110_SLICE_X21Y110_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_R_X15Y101_SLICE_X20Y101_AO6),
.I5(LIOB33_X0Y151_IOB_X0Y152_I),
.O5(CLBLM_R_X15Y110_SLICE_X20Y110_DO5),
.O6(CLBLM_R_X15Y110_SLICE_X20Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X15Y110_SLICE_X20Y110_CLUT (
.I0(CLBLM_R_X15Y110_SLICE_X20Y110_AO6),
.I1(CLBLM_R_X15Y109_SLICE_X20Y109_AO6),
.I2(CLBLM_R_X15Y109_SLICE_X20Y109_AO5),
.I3(CLBLM_R_X13Y109_SLICE_X18Y109_DO6),
.I4(CLBLM_R_X13Y113_SLICE_X19Y113_DO6),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_AO6),
.O5(CLBLM_R_X15Y110_SLICE_X20Y110_CO5),
.O6(CLBLM_R_X15Y110_SLICE_X20Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010005)
  ) CLBLM_R_X15Y110_SLICE_X20Y110_BLUT (
.I0(LIOB33_X0Y85_IOB_X0Y86_I),
.I1(LIOB33_X0Y65_IOB_X0Y66_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I4(LIOB33_X0Y71_IOB_X0Y71_I),
.I5(CLBLM_R_X15Y111_SLICE_X20Y111_AO6),
.O5(CLBLM_R_X15Y110_SLICE_X20Y110_BO5),
.O6(CLBLM_R_X15Y110_SLICE_X20Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h333301010000fafa)
  ) CLBLM_R_X15Y110_SLICE_X20Y110_ALUT (
.I0(LIOB33_X0Y87_IOB_X0Y88_I),
.I1(LIOB33_X0Y123_IOB_X0Y123_I),
.I2(LIOB33_X0Y89_IOB_X0Y90_I),
.I3(1'b1),
.I4(LIOB33_X0Y95_IOB_X0Y95_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y110_SLICE_X20Y110_AO5),
.O6(CLBLM_R_X15Y110_SLICE_X20Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff30ff0100000000)
  ) CLBLM_R_X15Y110_SLICE_X21Y110_DLUT (
.I0(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.I1(CLBLM_R_X13Y109_SLICE_X18Y109_DO6),
.I2(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.I3(CLBLM_R_X15Y111_SLICE_X21Y111_AO6),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O5(CLBLM_R_X15Y110_SLICE_X21Y110_DO5),
.O6(CLBLM_R_X15Y110_SLICE_X21Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0cc04cc00cc00)
  ) CLBLM_R_X15Y110_SLICE_X21Y110_CLUT (
.I0(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.I3(CLBLM_R_X15Y110_SLICE_X21Y110_AO5),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(CLBLM_R_X15Y99_SLICE_X20Y99_AO5),
.O5(CLBLM_R_X15Y110_SLICE_X21Y110_CO5),
.O6(CLBLM_R_X15Y110_SLICE_X21Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000076ff0000)
  ) CLBLM_R_X15Y110_SLICE_X21Y110_BLUT (
.I0(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.I1(LIOB33_X0Y125_IOB_X0Y126_I),
.I2(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.I3(CLBLM_R_X15Y99_SLICE_X20Y99_AO5),
.I4(CLBLM_R_X15Y110_SLICE_X21Y110_AO6),
.I5(RIOB33_X105Y167_IOB_X1Y167_I),
.O5(CLBLM_R_X15Y110_SLICE_X21Y110_BO5),
.O6(CLBLM_R_X15Y110_SLICE_X21Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f0f0ffffafafa)
  ) CLBLM_R_X15Y110_SLICE_X21Y110_ALUT (
.I0(RIOB33_X105Y167_IOB_X1Y167_I),
.I1(1'b1),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(LIOB33_X0Y65_IOB_X0Y66_I),
.I4(LIOB33_X0Y71_IOB_X0Y71_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y110_SLICE_X21Y110_AO5),
.O6(CLBLM_R_X15Y110_SLICE_X21Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y111_SLICE_X20Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y111_SLICE_X20Y111_DO5),
.O6(CLBLM_R_X15Y111_SLICE_X20Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y111_SLICE_X20Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y111_SLICE_X20Y111_CO5),
.O6(CLBLM_R_X15Y111_SLICE_X20Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0c0ccccc0c8c)
  ) CLBLM_R_X15Y111_SLICE_X20Y111_BLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(CLBLM_R_X15Y109_SLICE_X20Y109_AO6),
.I3(LIOB33_X0Y93_IOB_X0Y93_I),
.I4(LIOB33_X0Y127_IOB_X0Y128_I),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.O5(CLBLM_R_X15Y111_SLICE_X20Y111_BO5),
.O6(CLBLM_R_X15Y111_SLICE_X20Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff8ffffffffff)
  ) CLBLM_R_X15Y111_SLICE_X20Y111_ALUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(LIOB33_X0Y69_IOB_X0Y70_I),
.I2(LIOB33_X0Y91_IOB_X0Y91_I),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(LIOB33_X0Y87_IOB_X0Y88_I),
.I5(LIOB33_X0Y123_IOB_X0Y123_I),
.O5(CLBLM_R_X15Y111_SLICE_X20Y111_AO5),
.O6(CLBLM_R_X15Y111_SLICE_X20Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y111_SLICE_X21Y111_DO5),
.O6(CLBLM_R_X15Y111_SLICE_X21Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y111_SLICE_X21Y111_CO5),
.O6(CLBLM_R_X15Y111_SLICE_X21Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55557777fafafbfb)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_BLUT (
.I0(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.I1(LIOB33_X0Y123_IOB_X0Y123_I),
.I2(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.I3(1'b1),
.I4(CLBLM_R_X15Y110_SLICE_X20Y110_AO5),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLM_R_X15Y111_SLICE_X21Y111_BO5),
.O6(CLBLM_R_X15Y111_SLICE_X21Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff070700770077)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_ALUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(LIOB33_X0Y69_IOB_X0Y70_I),
.I2(LIOB33_X0Y85_IOB_X0Y86_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y165_IOB_X1Y165_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y111_SLICE_X21Y111_AO5),
.O6(CLBLM_R_X15Y111_SLICE_X21Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0202aaaa02aa)
  ) CLBLM_R_X15Y113_SLICE_X20Y113_DLUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I4(RIOB33_X105Y157_IOB_X1Y158_I),
.I5(CLBLM_R_X15Y113_SLICE_X20Y113_BO6),
.O5(CLBLM_R_X15Y113_SLICE_X20Y113_DO5),
.O6(CLBLM_R_X15Y113_SLICE_X20Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000fb000000f3)
  ) CLBLM_R_X15Y113_SLICE_X20Y113_CLUT (
.I0(LIOB33_X0Y151_IOB_X0Y151_I),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_DO6),
.I2(RIOB33_X105Y171_IOB_X1Y172_I),
.I3(LIOB33_X0Y159_IOB_X0Y160_I),
.I4(LIOB33_X0Y159_IOB_X0Y159_I),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLM_R_X15Y113_SLICE_X20Y113_CO5),
.O6(CLBLM_R_X15Y113_SLICE_X20Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafffff5f4f0f0)
  ) CLBLM_R_X15Y113_SLICE_X20Y113_BLUT (
.I0(LIOB33_X0Y55_IOB_X0Y56_I),
.I1(LIOB33_X0Y151_IOB_X0Y151_I),
.I2(RIOB33_X105Y157_IOB_X1Y158_I),
.I3(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X20Y113_BO5),
.O6(CLBLM_R_X15Y113_SLICE_X20Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffee0000cc88)
  ) CLBLM_R_X15Y113_SLICE_X20Y113_ALUT (
.I0(LIOB33_X0Y91_IOB_X0Y92_I),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(1'b1),
.I3(LIOB33_X0Y91_IOB_X0Y91_I),
.I4(LIOB33_X0Y95_IOB_X0Y95_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X20Y113_AO5),
.O6(CLBLM_R_X15Y113_SLICE_X20Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0c0f010)
  ) CLBLM_R_X15Y113_SLICE_X21Y113_DLUT (
.I0(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.I1(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I3(CLBLM_R_X15Y113_SLICE_X21Y113_AO5),
.I4(LIOB33_X0Y125_IOB_X0Y126_I),
.I5(CLBLM_R_X15Y113_SLICE_X20Y113_AO6),
.O5(CLBLM_R_X15Y113_SLICE_X21Y113_DO5),
.O6(CLBLM_R_X15Y113_SLICE_X21Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff000700)
  ) CLBLM_R_X15Y113_SLICE_X21Y113_CLUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(CLBLM_R_X13Y111_SLICE_X19Y111_AO5),
.I2(CLBLM_R_X15Y111_SLICE_X21Y111_BO6),
.I3(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I4(RIOB33_X105Y159_IOB_X1Y160_I),
.I5(CLBLM_R_X15Y113_SLICE_X21Y113_BO6),
.O5(CLBLM_R_X15Y113_SLICE_X21Y113_CO5),
.O6(CLBLM_R_X15Y113_SLICE_X21Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00007700f0f0f7f0)
  ) CLBLM_R_X15Y113_SLICE_X21Y113_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(LIOB33_X0Y69_IOB_X0Y70_I),
.I2(RIOB33_X105Y159_IOB_X1Y160_I),
.I3(LIOB33_X0Y123_IOB_X0Y123_I),
.I4(LIOB33_X0Y87_IOB_X0Y88_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X21Y113_BO5),
.O6(CLBLM_R_X15Y113_SLICE_X21Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888f0f0f7f0)
  ) CLBLM_R_X15Y113_SLICE_X21Y113_ALUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(LIOB33_X0Y69_IOB_X0Y70_I),
.I2(RIOB33_X105Y155_IOB_X1Y156_I),
.I3(LIOB33_X0Y125_IOB_X0Y125_I),
.I4(LIOB33_X0Y91_IOB_X0Y91_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X21Y113_AO5),
.O6(CLBLM_R_X15Y113_SLICE_X21Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505050004)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_DLUT (
.I0(LIOB33_X0Y159_IOB_X0Y160_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(LIOB33_X0Y159_IOB_X0Y159_I),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I4(RIOB33_X105Y157_IOB_X1Y157_I),
.I5(CLBLM_R_X15Y114_SLICE_X20Y114_BO6),
.O5(CLBLM_R_X15Y114_SLICE_X20Y114_DO5),
.O6(CLBLM_R_X15Y114_SLICE_X20Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000032323233)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_CLUT (
.I0(CLBLM_R_X15Y114_SLICE_X20Y114_AO6),
.I1(LIOB33_X0Y159_IOB_X0Y159_I),
.I2(RIOB33_X105Y159_IOB_X1Y159_I),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I5(LIOB33_X0Y159_IOB_X0Y160_I),
.O5(CLBLM_R_X15Y114_SLICE_X20Y114_CO5),
.O6(CLBLM_R_X15Y114_SLICE_X20Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030300045454555)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_BLUT (
.I0(RIOB33_X105Y157_IOB_X1Y157_I),
.I1(LIOB33_X0Y59_IOB_X0Y60_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y114_SLICE_X20Y114_BO5),
.O6(CLBLM_R_X15Y114_SLICE_X20Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a0a0a0ccececec)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(RIOB33_X105Y159_IOB_X1Y159_I),
.I2(LIOB33_X0Y119_IOB_X0Y119_I),
.I3(LIOB33_X0Y67_IOB_X0Y68_I),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(1'b1),
.O5(CLBLM_R_X15Y114_SLICE_X20Y114_AO5),
.O6(CLBLM_R_X15Y114_SLICE_X20Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y114_SLICE_X21Y114_DO5),
.O6(CLBLM_R_X15Y114_SLICE_X21Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y114_SLICE_X21Y114_CO5),
.O6(CLBLM_R_X15Y114_SLICE_X21Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y114_SLICE_X21Y114_BO5),
.O6(CLBLM_R_X15Y114_SLICE_X21Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y114_SLICE_X21Y114_AO5),
.O6(CLBLM_R_X15Y114_SLICE_X21Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X20Y123_DO5),
.O6(CLBLM_R_X15Y123_SLICE_X20Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X20Y123_CO5),
.O6(CLBLM_R_X15Y123_SLICE_X20Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X20Y123_BO5),
.O6(CLBLM_R_X15Y123_SLICE_X20Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f000f000f)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y159_IOB_X0Y160_I),
.I3(LIOB33_X0Y159_IOB_X0Y159_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X20Y123_AO5),
.O6(CLBLM_R_X15Y123_SLICE_X20Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X21Y123_DO5),
.O6(CLBLM_R_X15Y123_SLICE_X21Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X21Y123_CO5),
.O6(CLBLM_R_X15Y123_SLICE_X21Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X21Y123_BO5),
.O6(CLBLM_R_X15Y123_SLICE_X21Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X21Y123_AO5),
.O6(CLBLM_R_X15Y123_SLICE_X21Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300003332)
  ) CLBLM_R_X37Y111_SLICE_X56Y111_DLUT (
.I0(LIOB33_X0Y165_IOB_X0Y166_I),
.I1(LIOB33_X0Y157_IOB_X0Y158_I),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(CLBLM_R_X15Y113_SLICE_X20Y113_CO6),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.O5(CLBLM_R_X37Y111_SLICE_X56Y111_DO5),
.O6(CLBLM_R_X37Y111_SLICE_X56Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f00000f0e)
  ) CLBLM_R_X37Y111_SLICE_X56Y111_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y157_IOB_X0Y158_I),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(CLBLM_R_X15Y111_SLICE_X20Y111_BO6),
.O5(CLBLM_R_X37Y111_SLICE_X56Y111_CO5),
.O6(CLBLM_R_X37Y111_SLICE_X56Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff00fe)
  ) CLBLM_R_X37Y111_SLICE_X56Y111_BLUT (
.I0(LIOB33_X0Y51_IOB_X0Y51_I),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I2(CLBLM_R_X15Y113_SLICE_X20Y113_CO6),
.I3(LIOB33_X0Y153_IOB_X0Y154_I),
.I4(LIOB33_X0Y165_IOB_X0Y166_I),
.I5(LIOB33_X0Y155_IOB_X0Y156_I),
.O5(CLBLM_R_X37Y111_SLICE_X56Y111_BO5),
.O6(CLBLM_R_X37Y111_SLICE_X56Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500550054)
  ) CLBLM_R_X37Y111_SLICE_X56Y111_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_R_X15Y111_SLICE_X20Y111_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y155_IOB_X0Y156_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.O5(CLBLM_R_X37Y111_SLICE_X56Y111_AO5),
.O6(CLBLM_R_X37Y111_SLICE_X56Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y111_SLICE_X57Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y111_SLICE_X57Y111_DO5),
.O6(CLBLM_R_X37Y111_SLICE_X57Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y111_SLICE_X57Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y111_SLICE_X57Y111_CO5),
.O6(CLBLM_R_X37Y111_SLICE_X57Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y111_SLICE_X57Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y111_SLICE_X57Y111_BO5),
.O6(CLBLM_R_X37Y111_SLICE_X57Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y111_SLICE_X57Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y111_SLICE_X57Y111_AO5),
.O6(CLBLM_R_X37Y111_SLICE_X57Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X146Y116_DO5),
.O6(CLBLM_R_X93Y116_SLICE_X146Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X146Y116_CO5),
.O6(CLBLM_R_X93Y116_SLICE_X146Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X146Y116_BO5),
.O6(CLBLM_R_X93Y116_SLICE_X146Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X146Y116_AO5),
.O6(CLBLM_R_X93Y116_SLICE_X146Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X147Y116_DO5),
.O6(CLBLM_R_X93Y116_SLICE_X147Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X147Y116_CO5),
.O6(CLBLM_R_X93Y116_SLICE_X147Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X147Y116_BO5),
.O6(CLBLM_R_X93Y116_SLICE_X147Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefcfcfefffcfc)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_ALUT (
.I0(CLBLM_R_X15Y113_SLICE_X21Y113_BO5),
.I1(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(CLBLM_R_X15Y111_SLICE_X21Y111_BO6),
.I4(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I5(CLBLM_R_X15Y113_SLICE_X20Y113_AO5),
.O5(CLBLM_R_X93Y116_SLICE_X147Y116_AO5),
.O6(CLBLM_R_X93Y116_SLICE_X147Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X146Y122_DO5),
.O6(CLBLM_R_X93Y122_SLICE_X146Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X146Y122_CO5),
.O6(CLBLM_R_X93Y122_SLICE_X146Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X146Y122_BO5),
.O6(CLBLM_R_X93Y122_SLICE_X146Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X146Y122_AO5),
.O6(CLBLM_R_X93Y122_SLICE_X146Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X147Y122_DO5),
.O6(CLBLM_R_X93Y122_SLICE_X147Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccc040000)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I1(CLBLL_R_X81Y122_SLICE_X126Y122_CO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I4(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I5(CLBLM_R_X93Y122_SLICE_X147Y122_BO6),
.O5(CLBLM_R_X93Y122_SLICE_X147Y122_CO5),
.O6(CLBLM_R_X93Y122_SLICE_X147Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffccffefffcc)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_BLUT (
.I0(CLBLM_R_X15Y113_SLICE_X21Y113_BO5),
.I1(RIOB33_X105Y151_IOB_X1Y151_I),
.I2(CLBLM_R_X15Y111_SLICE_X21Y111_BO6),
.I3(RIOB33_X105Y151_IOB_X1Y152_I),
.I4(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I5(CLBLM_R_X15Y113_SLICE_X20Y113_AO5),
.O5(CLBLM_R_X93Y122_SLICE_X147Y122_BO5),
.O6(CLBLM_R_X93Y122_SLICE_X147Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa0000ff020000)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_ALUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I3(CLBLM_R_X93Y122_SLICE_X147Y122_BO6),
.I4(CLBLL_R_X81Y124_SLICE_X126Y124_AO6),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O5(CLBLM_R_X93Y122_SLICE_X147Y122_AO5),
.O6(CLBLM_R_X93Y122_SLICE_X147Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_DO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_CO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_BO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefefeffffffaa)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_ALUT (
.I0(CLBLM_R_X15Y110_SLICE_X21Y110_DO6),
.I1(LIOB33_X0Y121_IOB_X0Y121_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(RIOB33_X105Y125_IOB_X1Y126_I),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_AO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_DO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_CO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_BO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_AO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e0c0c0e0e0c0e0)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_DLUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I1(CLBLM_R_X101Y123_SLICE_X158Y123_AO5),
.I2(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I4(CLBLM_R_X15Y113_SLICE_X20Y113_BO5),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.O5(CLBLM_R_X101Y124_SLICE_X158Y124_DO5),
.O6(CLBLM_R_X101Y124_SLICE_X158Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hecec0000ecee0000)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_CLUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I1(CLBLM_R_X101Y123_SLICE_X158Y123_AO5),
.I2(CLBLM_R_X15Y113_SLICE_X20Y113_BO5),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I4(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.O5(CLBLM_R_X101Y124_SLICE_X158Y124_CO5),
.O6(CLBLM_R_X101Y124_SLICE_X158Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a000ff00b000)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_BLUT (
.I0(CLBLM_R_X15Y113_SLICE_X20Y113_BO5),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I3(CLBLL_R_X81Y122_SLICE_X126Y122_CO6),
.I4(CLBLM_R_X101Y123_SLICE_X158Y123_AO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O5(CLBLM_R_X101Y124_SLICE_X158Y124_BO5),
.O6(CLBLM_R_X101Y124_SLICE_X158Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f08080f0f080c0)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_ALUT (
.I0(CLBLM_R_X15Y113_SLICE_X20Y113_BO5),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I2(CLBLL_R_X81Y124_SLICE_X126Y124_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I4(CLBLM_R_X101Y123_SLICE_X158Y123_AO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O5(CLBLM_R_X101Y124_SLICE_X158Y124_AO5),
.O6(CLBLM_R_X101Y124_SLICE_X158Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X159Y124_DO5),
.O6(CLBLM_R_X101Y124_SLICE_X159Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X159Y124_CO5),
.O6(CLBLM_R_X101Y124_SLICE_X159Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X159Y124_BO5),
.O6(CLBLM_R_X101Y124_SLICE_X159Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X159Y124_AO5),
.O6(CLBLM_R_X101Y124_SLICE_X159Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X162Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X162Y97_DO5),
.O6(CLBLM_R_X103Y97_SLICE_X162Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X162Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X162Y97_CO5),
.O6(CLBLM_R_X103Y97_SLICE_X162Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X162Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X162Y97_BO5),
.O6(CLBLM_R_X103Y97_SLICE_X162Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X162Y97_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X162Y97_AO5),
.O6(CLBLM_R_X103Y97_SLICE_X162Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X163Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X163Y97_DO5),
.O6(CLBLM_R_X103Y97_SLICE_X163Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X163Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X163Y97_CO5),
.O6(CLBLM_R_X103Y97_SLICE_X163Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fe00fe00)
  ) CLBLM_R_X103Y97_SLICE_X163Y97_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I1(CLBLM_R_X15Y111_SLICE_X20Y111_BO6),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.I4(1'b1),
.I5(LIOB33_X0Y51_IOB_X0Y52_I),
.O5(CLBLM_R_X103Y97_SLICE_X163Y97_BO5),
.O6(CLBLM_R_X103Y97_SLICE_X163Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fe00fe00)
  ) CLBLM_R_X103Y97_SLICE_X163Y97_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I1(CLBLM_R_X15Y111_SLICE_X20Y111_BO6),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y51_IOB_X0Y52_I),
.O5(CLBLM_R_X103Y97_SLICE_X163Y97_AO5),
.O6(CLBLM_R_X103Y97_SLICE_X163Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y103_SLICE_X162Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y103_SLICE_X162Y103_DO5),
.O6(CLBLM_R_X103Y103_SLICE_X162Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y103_SLICE_X162Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y103_SLICE_X162Y103_CO5),
.O6(CLBLM_R_X103Y103_SLICE_X162Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y103_SLICE_X162Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y103_SLICE_X162Y103_BO5),
.O6(CLBLM_R_X103Y103_SLICE_X162Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y103_SLICE_X162Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y103_SLICE_X162Y103_AO5),
.O6(CLBLM_R_X103Y103_SLICE_X162Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y103_SLICE_X163Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y103_SLICE_X163Y103_DO5),
.O6(CLBLM_R_X103Y103_SLICE_X163Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y103_SLICE_X163Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y103_SLICE_X163Y103_CO5),
.O6(CLBLM_R_X103Y103_SLICE_X163Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaaaaa0)
  ) CLBLM_R_X103Y103_SLICE_X163Y103_BLUT (
.I0(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.I1(1'b1),
.I2(CLBLM_R_X15Y113_SLICE_X20Y113_CO6),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X103Y103_SLICE_X163Y103_BO5),
.O6(CLBLM_R_X103Y103_SLICE_X163Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffee0000)
  ) CLBLM_R_X103Y103_SLICE_X163Y103_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.I5(CLBLM_R_X15Y113_SLICE_X20Y113_CO6),
.O5(CLBLM_R_X103Y103_SLICE_X163Y103_AO5),
.O6(CLBLM_R_X103Y103_SLICE_X163Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X162Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X162Y107_DO5),
.O6(CLBLM_R_X103Y107_SLICE_X162Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X162Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X162Y107_CO5),
.O6(CLBLM_R_X103Y107_SLICE_X162Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X162Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X162Y107_BO5),
.O6(CLBLM_R_X103Y107_SLICE_X162Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X162Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X162Y107_AO5),
.O6(CLBLM_R_X103Y107_SLICE_X162Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X163Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X163Y107_DO5),
.O6(CLBLM_R_X103Y107_SLICE_X163Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X163Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X163Y107_CO5),
.O6(CLBLM_R_X103Y107_SLICE_X163Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfd00000000)
  ) CLBLM_R_X103Y107_SLICE_X163Y107_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_DO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(1'b1),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.O5(CLBLM_R_X103Y107_SLICE_X163Y107_BO5),
.O6(CLBLM_R_X103Y107_SLICE_X163Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fd0055555555)
  ) CLBLM_R_X103Y107_SLICE_X163Y107_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_DO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X163Y107_AO5),
.O6(CLBLM_R_X103Y107_SLICE_X163Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_DO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_CO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_BO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_AO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_DO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00ee00)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_CO6),
.I2(1'b1),
.I3(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.I4(RIOB33_X105Y123_IOB_X1Y124_I),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_CO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffe00000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_BLUT (
.I0(RIOB33_X105Y123_IOB_X1Y124_I),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLM_R_X13Y113_SLICE_X19Y113_CO6),
.I4(1'b1),
.I5(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_BO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cc00cc00)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(1'b1),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_AO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_DO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_CO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_BO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_AO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_DO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_CO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_ALUT (
.I0(RIOB33_X105Y123_IOB_X1Y123_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y121_IOB_X1Y122_I),
.I5(CLBLM_R_X13Y110_SLICE_X19Y110_CO6),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X162Y125_DO5),
.O6(CLBLM_R_X103Y125_SLICE_X162Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X162Y125_CO5),
.O6(CLBLM_R_X103Y125_SLICE_X162Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f8fa00000000)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_BLUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I1(CLBLM_R_X15Y114_SLICE_X20Y114_AO5),
.I2(CLBLM_R_X103Y125_SLICE_X163Y125_AO5),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I5(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.O5(CLBLM_R_X103Y125_SLICE_X162Y125_BO5),
.O6(CLBLM_R_X103Y125_SLICE_X162Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf080f080f080f0a0)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_ALUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.I1(CLBLM_R_X15Y114_SLICE_X20Y114_AO5),
.I2(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.I3(CLBLM_R_X103Y125_SLICE_X163Y125_AO5),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.O5(CLBLM_R_X103Y125_SLICE_X162Y125_AO5),
.O6(CLBLM_R_X103Y125_SLICE_X162Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X163Y125_DO5),
.O6(CLBLM_R_X103Y125_SLICE_X163Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X163Y125_CO5),
.O6(CLBLM_R_X103Y125_SLICE_X163Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X163Y125_BO5),
.O6(CLBLM_R_X103Y125_SLICE_X163Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefefeffffffaa)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_ALUT (
.I0(CLBLM_R_X15Y110_SLICE_X21Y110_CO6),
.I1(RIOB33_X105Y153_IOB_X1Y154_I),
.I2(RIOB33_X105Y153_IOB_X1Y153_I),
.I3(RIOB33_X105Y125_IOB_X1Y125_I),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X163Y125_AO5),
.O6(CLBLM_R_X103Y125_SLICE_X163Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X162Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X162Y147_DO5),
.O6(CLBLM_R_X103Y147_SLICE_X162Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X162Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X162Y147_CO5),
.O6(CLBLM_R_X103Y147_SLICE_X162Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X162Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X162Y147_BO5),
.O6(CLBLM_R_X103Y147_SLICE_X162Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X162Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X162Y147_AO5),
.O6(CLBLM_R_X103Y147_SLICE_X162Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X163Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X163Y147_DO5),
.O6(CLBLM_R_X103Y147_SLICE_X163Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X163Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X163Y147_CO5),
.O6(CLBLM_R_X103Y147_SLICE_X163Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X163Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X163Y147_BO5),
.O6(CLBLM_R_X103Y147_SLICE_X163Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888833333333)
  ) CLBLM_R_X103Y147_SLICE_X163Y147_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y147_IOB_X0Y147_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X163Y147_AO5),
.O6(CLBLM_R_X103Y147_SLICE_X163Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f55555555)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(RIOB33_SING_X105Y150_IOB_X1Y150_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X162Y185_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X162Y185_DO5),
.O6(CLBLM_R_X103Y185_SLICE_X162Y185_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X162Y185_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X162Y185_CO5),
.O6(CLBLM_R_X103Y185_SLICE_X162Y185_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X162Y185_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X162Y185_BO5),
.O6(CLBLM_R_X103Y185_SLICE_X162Y185_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X162Y185_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X162Y185_AO5),
.O6(CLBLM_R_X103Y185_SLICE_X162Y185_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X163Y185_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X163Y185_DO5),
.O6(CLBLM_R_X103Y185_SLICE_X163Y185_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X163Y185_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X163Y185_CO5),
.O6(CLBLM_R_X103Y185_SLICE_X163Y185_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X163Y185_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X163Y185_BO5),
.O6(CLBLM_R_X103Y185_SLICE_X163Y185_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X103Y185_SLICE_X163Y185_ALUT (
.I0(LIOB33_X0Y133_IOB_X0Y134_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X163Y185_AO5),
.O6(CLBLM_R_X103Y185_SLICE_X163Y185_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y80_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y80_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y81_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y81_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y82_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y82_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y82_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y83_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y83_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y83_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y84_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y84_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y84_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y85_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y85_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y86_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y86_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y86_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y87_IOB_X0Y87_IBUF (
.I(LIOB33_X0Y87_IOB_X0Y87_IPAD),
.O(LIOB33_X0Y87_IOB_X0Y87_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y87_IOB_X0Y88_IBUF (
.I(LIOB33_X0Y87_IOB_X0Y88_IPAD),
.O(LIOB33_X0Y87_IOB_X0Y88_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y89_IOB_X0Y89_IBUF (
.I(LIOB33_X0Y89_IOB_X0Y89_IPAD),
.O(LIOB33_X0Y89_IOB_X0Y89_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y89_IOB_X0Y90_IBUF (
.I(LIOB33_X0Y89_IOB_X0Y90_IPAD),
.O(LIOB33_X0Y89_IOB_X0Y90_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y91_IOB_X0Y91_IBUF (
.I(LIOB33_X0Y91_IOB_X0Y91_IPAD),
.O(LIOB33_X0Y91_IOB_X0Y91_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y91_IOB_X0Y92_IBUF (
.I(LIOB33_X0Y91_IOB_X0Y92_IPAD),
.O(LIOB33_X0Y91_IOB_X0Y92_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y93_IOB_X0Y93_IBUF (
.I(LIOB33_X0Y93_IOB_X0Y93_IPAD),
.O(LIOB33_X0Y93_IOB_X0Y93_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y93_IOB_X0Y94_IBUF (
.I(LIOB33_X0Y93_IOB_X0Y94_IPAD),
.O(LIOB33_X0Y93_IOB_X0Y94_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y95_IOB_X0Y95_IBUF (
.I(LIOB33_X0Y95_IOB_X0Y95_IPAD),
.O(LIOB33_X0Y95_IOB_X0Y95_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y95_IOB_X0Y96_IBUF (
.I(LIOB33_X0Y95_IOB_X0Y96_IPAD),
.O(LIOB33_X0Y95_IOB_X0Y96_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y97_IOB_X0Y97_IBUF (
.I(LIOB33_X0Y97_IOB_X0Y97_IPAD),
.O(LIOB33_X0Y97_IOB_X0Y97_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y97_IOB_X0Y98_IBUF (
.I(LIOB33_X0Y97_IOB_X0Y98_IPAD),
.O(LIOB33_X0Y97_IOB_X0Y98_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y124_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y126_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y127_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y129_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y129_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y130_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y130_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y131_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y131_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y132_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y132_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y133_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y134_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y135_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y136_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y136_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(LIOB33_X0Y137_IOB_X0Y137_IPAD),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y137_IOB_X0Y138_IBUF (
.I(LIOB33_X0Y137_IOB_X0Y138_IPAD),
.O(LIOB33_X0Y137_IOB_X0Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y139_IOB_X0Y139_IBUF (
.I(LIOB33_X0Y139_IOB_X0Y139_IPAD),
.O(LIOB33_X0Y139_IOB_X0Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y139_IOB_X0Y140_IBUF (
.I(LIOB33_X0Y139_IOB_X0Y140_IPAD),
.O(LIOB33_X0Y139_IOB_X0Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y141_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y141_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y142_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y142_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y143_IOB_X0Y143_IBUF (
.I(LIOB33_X0Y143_IOB_X0Y143_IPAD),
.O(LIOB33_X0Y143_IOB_X0Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y145_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y145_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y146_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y146_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y147_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y147_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y148_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y148_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y151_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y151_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y152_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y152_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y153_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y153_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y154_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y154_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y155_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y156_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y156_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y157_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y157_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y158_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y158_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y159_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y159_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y160_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y160_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y161_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y161_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y162_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y162_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y163_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y163_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y164_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y164_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y165_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y165_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y166_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y166_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y167_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y167_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y168_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y168_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y169_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y169_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y170_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y170_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y171_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y171_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y172_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y172_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y173_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y173_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y173_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y174_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y174_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y174_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y175_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y175_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y175_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y176_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y176_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y176_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y177_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y177_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y177_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(CLBLL_L_X2Y175_SLICE_X0Y175_AO6),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(LIOB33_X0Y97_IOB_X0Y97_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(CLBLM_R_X103Y108_SLICE_X163Y108_AO5),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(CLBLL_L_X2Y174_SLICE_X0Y174_BO6),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(CLBLL_L_X2Y174_SLICE_X0Y174_BO6),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(CLBLL_L_X2Y174_SLICE_X0Y174_BO6),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(CLBLL_L_X2Y174_SLICE_X0Y174_BO6),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(1'b0),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(1'b0),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(CLBLL_L_X2Y101_SLICE_X0Y101_BO6),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y99_IOB_X0Y99_IBUF (
.I(LIOB33_SING_X0Y99_IOB_X0Y99_IPAD),
.O(LIOB33_SING_X0Y99_IOB_X0Y99_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y149_IOB_X0Y149_IBUF (
.I(LIOB33_SING_X0Y149_IOB_X0Y149_IPAD),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y150_IOB_X0Y150_IBUF (
.I(LIOB33_SING_X0Y150_IOB_X0Y150_IPAD),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y200_IOB_X0Y200_OBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O(LIOB33_SING_X0Y200_IOB_X0Y200_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y51_OBUF (
.I(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.O(RIOB33_X105Y51_IOB_X1Y51_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y52_OBUF (
.I(CLBLM_R_X15Y99_SLICE_X20Y99_AO6),
.O(RIOB33_X105Y51_IOB_X1Y52_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y53_OBUF (
.I(CLBLM_R_X13Y110_SLICE_X19Y110_CO6),
.O(RIOB33_X105Y53_IOB_X1Y53_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y54_OBUF (
.I(CLBLM_R_X103Y108_SLICE_X163Y108_AO6),
.O(RIOB33_X105Y53_IOB_X1Y54_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y55_OBUF (
.I(CLBLM_R_X13Y113_SLICE_X19Y113_CO6),
.O(RIOB33_X105Y55_IOB_X1Y55_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y56_OBUF (
.I(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.O(RIOB33_X105Y55_IOB_X1Y56_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y57_OBUF (
.I(CLBLM_R_X15Y109_SLICE_X20Y109_BO6),
.O(RIOB33_X105Y57_IOB_X1Y57_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y58_OBUF (
.I(CLBLL_R_X81Y122_SLICE_X126Y122_AO6),
.O(RIOB33_X105Y57_IOB_X1Y58_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y59_OBUF (
.I(CLBLM_R_X15Y111_SLICE_X20Y111_BO6),
.O(RIOB33_X105Y59_IOB_X1Y59_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y60_OBUF (
.I(CLBLM_R_X15Y113_SLICE_X20Y113_CO6),
.O(RIOB33_X105Y59_IOB_X1Y60_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y61_OBUF (
.I(CLBLM_R_X13Y112_SLICE_X19Y112_DO6),
.O(RIOB33_X105Y61_IOB_X1Y61_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y62_OBUF (
.I(CLBLL_R_X81Y122_SLICE_X126Y122_BO6),
.O(RIOB33_X105Y61_IOB_X1Y62_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y63_OBUF (
.I(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.O(RIOB33_X105Y63_IOB_X1Y63_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y64_OBUF (
.I(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.O(RIOB33_X105Y63_IOB_X1Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y65_OBUF (
.I(CLBLM_R_X103Y107_SLICE_X163Y107_AO5),
.O(RIOB33_X105Y65_IOB_X1Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y66_OBUF (
.I(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.O(RIOB33_X105Y65_IOB_X1Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y67_OBUF (
.I(CLBLM_R_X13Y109_SLICE_X18Y109_AO6),
.O(RIOB33_X105Y67_IOB_X1Y67_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y68_OBUF (
.I(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.O(RIOB33_X105Y67_IOB_X1Y68_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y69_OBUF (
.I(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.O(RIOB33_X105Y69_IOB_X1Y69_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y70_OBUF (
.I(CLBLM_R_X15Y110_SLICE_X20Y110_CO6),
.O(RIOB33_X105Y69_IOB_X1Y70_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y71_OBUF (
.I(CLBLM_L_X92Y125_SLICE_X144Y125_AO6),
.O(RIOB33_X105Y71_IOB_X1Y71_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y72_OBUF (
.I(CLBLM_L_X92Y125_SLICE_X144Y125_BO6),
.O(RIOB33_X105Y71_IOB_X1Y72_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y73_OBUF (
.I(CLBLM_R_X37Y111_SLICE_X56Y111_BO6),
.O(RIOB33_X105Y73_IOB_X1Y73_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y74_OBUF (
.I(CLBLL_R_X81Y111_SLICE_X126Y111_AO6),
.O(RIOB33_X105Y73_IOB_X1Y74_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y75_OBUF (
.I(CLBLM_L_X30Y111_SLICE_X44Y111_AO6),
.O(RIOB33_X105Y75_IOB_X1Y75_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y76_OBUF (
.I(CLBLM_R_X37Y111_SLICE_X56Y111_CO6),
.O(RIOB33_X105Y75_IOB_X1Y76_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y77_OBUF (
.I(CLBLM_R_X37Y111_SLICE_X56Y111_DO6),
.O(RIOB33_X105Y77_IOB_X1Y77_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y78_OBUF (
.I(CLBLL_R_X81Y111_SLICE_X126Y111_BO6),
.O(RIOB33_X105Y77_IOB_X1Y78_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y79_OBUF (
.I(CLBLM_L_X30Y111_SLICE_X44Y111_BO6),
.O(RIOB33_X105Y79_IOB_X1Y79_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y80_OBUF (
.I(CLBLM_R_X103Y97_SLICE_X163Y97_AO6),
.O(RIOB33_X105Y79_IOB_X1Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y81_OBUF (
.I(CLBLM_R_X103Y108_SLICE_X163Y108_BO6),
.O(RIOB33_X105Y81_IOB_X1Y81_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y82_OBUF (
.I(CLBLM_R_X103Y107_SLICE_X163Y107_BO6),
.O(RIOB33_X105Y81_IOB_X1Y82_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y83_OBUF (
.I(CLBLM_R_X103Y103_SLICE_X163Y103_AO6),
.O(RIOB33_X105Y83_IOB_X1Y83_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y84_OBUF (
.I(CLBLM_R_X103Y97_SLICE_X163Y97_BO6),
.O(RIOB33_X105Y83_IOB_X1Y84_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y85_OBUF (
.I(CLBLM_R_X103Y108_SLICE_X163Y108_CO6),
.O(RIOB33_X105Y85_IOB_X1Y85_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y86_OBUF (
.I(CLBLM_R_X103Y107_SLICE_X163Y107_AO6),
.O(RIOB33_X105Y85_IOB_X1Y86_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y87_OBUF (
.I(CLBLM_R_X103Y103_SLICE_X163Y103_BO6),
.O(RIOB33_X105Y87_IOB_X1Y87_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y88_OBUF (
.I(CLBLM_R_X15Y110_SLICE_X20Y110_DO6),
.O(RIOB33_X105Y87_IOB_X1Y88_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y89_OBUF (
.I(CLBLM_R_X15Y101_SLICE_X20Y101_AO5),
.O(RIOB33_X105Y89_IOB_X1Y89_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y90_OBUF (
.I(CLBLM_R_X15Y110_SLICE_X21Y110_CO6),
.O(RIOB33_X105Y89_IOB_X1Y90_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y91_OBUF (
.I(CLBLM_R_X15Y110_SLICE_X21Y110_DO6),
.O(RIOB33_X105Y91_IOB_X1Y91_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y92_OBUF (
.I(CLBLM_R_X15Y113_SLICE_X21Y113_CO6),
.O(RIOB33_X105Y91_IOB_X1Y92_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y93_OBUF (
.I(CLBLM_R_X15Y113_SLICE_X21Y113_DO6),
.O(RIOB33_X105Y93_IOB_X1Y93_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y94_OBUF (
.I(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O(RIOB33_X105Y93_IOB_X1Y94_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y95_OBUF (
.I(CLBLM_R_X15Y114_SLICE_X20Y114_CO6),
.O(RIOB33_X105Y95_IOB_X1Y95_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y96_OBUF (
.I(CLBLM_R_X15Y113_SLICE_X20Y113_DO6),
.O(RIOB33_X105Y95_IOB_X1Y96_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y97_OBUF (
.I(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.O(RIOB33_X105Y97_IOB_X1Y97_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y98_OBUF (
.I(CLBLM_R_X15Y114_SLICE_X20Y114_DO6),
.O(RIOB33_X105Y97_IOB_X1Y98_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLM_R_X37Y111_SLICE_X56Y111_AO6),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y128_OBUF (
.I(CLBLL_L_X102Y125_SLICE_X161Y125_AO6),
.O(RIOB33_X105Y127_IOB_X1Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLL_L_X102Y125_SLICE_X161Y125_BO6),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLM_R_X101Y124_SLICE_X158Y124_AO6),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLM_R_X93Y122_SLICE_X147Y122_AO6),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLM_L_X78Y119_SLICE_X121Y119_AO6),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_R_X101Y124_SLICE_X158Y124_BO6),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLM_R_X93Y122_SLICE_X147Y122_CO6),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLM_L_X78Y119_SLICE_X121Y119_CO6),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(CLBLM_L_X94Y122_SLICE_X148Y122_AO6),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(CLBLM_R_X101Y124_SLICE_X158Y124_CO6),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(CLBLM_R_X103Y125_SLICE_X162Y125_AO6),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(CLBLM_L_X78Y119_SLICE_X121Y119_DO6),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLM_L_X94Y122_SLICE_X148Y122_BO6),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLM_R_X101Y124_SLICE_X158Y124_DO6),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLM_R_X103Y125_SLICE_X162Y125_BO6),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLM_L_X78Y125_SLICE_X121Y125_AO6),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(CLBLM_L_X78Y125_SLICE_X121Y125_BO6),
.O(RIOB33_X105Y145_IOB_X1Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLM_L_X78Y125_SLICE_X121Y125_CO6),
.O(RIOB33_X105Y147_IOB_X1Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLM_L_X78Y125_SLICE_X121Y125_DO6),
.O(RIOB33_X105Y147_IOB_X1Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y151_IOB_X1Y151_IBUF (
.I(RIOB33_X105Y151_IOB_X1Y151_IPAD),
.O(RIOB33_X105Y151_IOB_X1Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y151_IOB_X1Y152_IBUF (
.I(RIOB33_X105Y151_IOB_X1Y152_IPAD),
.O(RIOB33_X105Y151_IOB_X1Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y153_IOB_X1Y153_IBUF (
.I(RIOB33_X105Y153_IOB_X1Y153_IPAD),
.O(RIOB33_X105Y153_IOB_X1Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y153_IOB_X1Y154_IBUF (
.I(RIOB33_X105Y153_IOB_X1Y154_IPAD),
.O(RIOB33_X105Y153_IOB_X1Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y155_IOB_X1Y155_IBUF (
.I(RIOB33_X105Y155_IOB_X1Y155_IPAD),
.O(RIOB33_X105Y155_IOB_X1Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y155_IOB_X1Y156_IBUF (
.I(RIOB33_X105Y155_IOB_X1Y156_IPAD),
.O(RIOB33_X105Y155_IOB_X1Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y157_IOB_X1Y157_IBUF (
.I(RIOB33_X105Y157_IOB_X1Y157_IPAD),
.O(RIOB33_X105Y157_IOB_X1Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y157_IOB_X1Y158_IBUF (
.I(RIOB33_X105Y157_IOB_X1Y158_IPAD),
.O(RIOB33_X105Y157_IOB_X1Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y159_IOB_X1Y159_IBUF (
.I(RIOB33_X105Y159_IOB_X1Y159_IPAD),
.O(RIOB33_X105Y159_IOB_X1Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y159_IOB_X1Y160_IBUF (
.I(RIOB33_X105Y159_IOB_X1Y160_IPAD),
.O(RIOB33_X105Y159_IOB_X1Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y161_IOB_X1Y161_IBUF (
.I(RIOB33_X105Y161_IOB_X1Y161_IPAD),
.O(RIOB33_X105Y161_IOB_X1Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y161_IOB_X1Y162_IBUF (
.I(RIOB33_X105Y161_IOB_X1Y162_IPAD),
.O(RIOB33_X105Y161_IOB_X1Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y163_IOB_X1Y163_IBUF (
.I(RIOB33_X105Y163_IOB_X1Y163_IPAD),
.O(RIOB33_X105Y163_IOB_X1Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y163_IOB_X1Y164_IBUF (
.I(RIOB33_X105Y163_IOB_X1Y164_IPAD),
.O(RIOB33_X105Y163_IOB_X1Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y165_IOB_X1Y165_IBUF (
.I(RIOB33_X105Y165_IOB_X1Y165_IPAD),
.O(RIOB33_X105Y165_IOB_X1Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y165_IOB_X1Y166_IBUF (
.I(RIOB33_X105Y165_IOB_X1Y166_IPAD),
.O(RIOB33_X105Y165_IOB_X1Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y167_IOB_X1Y167_IBUF (
.I(RIOB33_X105Y167_IOB_X1Y167_IPAD),
.O(RIOB33_X105Y167_IOB_X1Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y167_IOB_X1Y168_IBUF (
.I(RIOB33_X105Y167_IOB_X1Y168_IPAD),
.O(RIOB33_X105Y167_IOB_X1Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y169_IOB_X1Y169_IBUF (
.I(RIOB33_X105Y169_IOB_X1Y169_IPAD),
.O(RIOB33_X105Y169_IOB_X1Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y169_IOB_X1Y170_IBUF (
.I(RIOB33_X105Y169_IOB_X1Y170_IPAD),
.O(RIOB33_X105Y169_IOB_X1Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y171_IOB_X1Y171_IBUF (
.I(RIOB33_X105Y171_IOB_X1Y171_IPAD),
.O(RIOB33_X105Y171_IOB_X1Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y171_IOB_X1Y172_IBUF (
.I(RIOB33_X105Y171_IOB_X1Y172_IPAD),
.O(RIOB33_X105Y171_IOB_X1Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y147_SLICE_X163Y147_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_I),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_I),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(LIOB33_X0Y137_IOB_X0Y138_I),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(LIOB33_X0Y137_IOB_X0Y137_I),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X103Y147_SLICE_X163Y147_AO6),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X0Y146_AO5),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLL_L_X2Y136_SLICE_X0Y136_BO6),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(RIOB33_SING_X105Y150_IOB_X1Y150_I),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_I),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_I),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X103Y185_SLICE_X163Y185_AO6),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X0Y146_AO6),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLL_L_X2Y174_SLICE_X0Y174_AO5),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X13Y110_SLICE_X19Y110_AO6),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_I),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X0Y173_AO6),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLL_L_X2Y174_SLICE_X0Y174_AO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLL_L_X2Y174_SLICE_X0Y174_AO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y50_IOB_X1Y50_OBUF (
.I(CLBLM_R_X15Y99_SLICE_X20Y99_AO6),
.O(RIOB33_SING_X105Y50_IOB_X1Y50_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y99_IOB_X1Y99_OBUF (
.I(CLBLM_L_X78Y119_SLICE_X121Y119_BO6),
.O(RIOB33_SING_X105Y99_IOB_X1Y99_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y150_IOB_X1Y150_IBUF (
.I(RIOB33_SING_X105Y150_IOB_X1Y150_IPAD),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLL_L_X2Y174_SLICE_X0Y174_BO5),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y101_SLICE_X0Y101_A = CLBLL_L_X2Y101_SLICE_X0Y101_AO6;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_B = CLBLL_L_X2Y101_SLICE_X0Y101_BO6;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_C = CLBLL_L_X2Y101_SLICE_X0Y101_CO6;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_D = CLBLL_L_X2Y101_SLICE_X0Y101_DO6;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_A = CLBLL_L_X2Y101_SLICE_X1Y101_AO6;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_B = CLBLL_L_X2Y101_SLICE_X1Y101_BO6;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_C = CLBLL_L_X2Y101_SLICE_X1Y101_CO6;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_D = CLBLL_L_X2Y101_SLICE_X1Y101_DO6;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A = CLBLL_L_X2Y136_SLICE_X0Y136_AO6;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B = CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C = CLBLL_L_X2Y136_SLICE_X0Y136_CO6;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D = CLBLL_L_X2Y136_SLICE_X0Y136_DO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A = CLBLL_L_X2Y136_SLICE_X1Y136_AO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B = CLBLL_L_X2Y136_SLICE_X1Y136_BO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C = CLBLL_L_X2Y136_SLICE_X1Y136_CO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D = CLBLL_L_X2Y136_SLICE_X1Y136_DO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B = CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C = CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D = CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_AMUX = CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A = CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B = CLBLL_L_X2Y173_SLICE_X0Y173_BO6;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C = CLBLL_L_X2Y173_SLICE_X0Y173_CO6;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D = CLBLL_L_X2Y173_SLICE_X0Y173_DO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A = CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C = CLBLL_L_X2Y173_SLICE_X1Y173_CO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D = CLBLL_L_X2Y173_SLICE_X1Y173_DO6;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_A = CLBLL_L_X2Y174_SLICE_X0Y174_AO6;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_B = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_C = CLBLL_L_X2Y174_SLICE_X0Y174_CO6;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_D = CLBLL_L_X2Y174_SLICE_X0Y174_DO6;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_AMUX = CLBLL_L_X2Y174_SLICE_X0Y174_AO5;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_BMUX = CLBLL_L_X2Y174_SLICE_X0Y174_BO5;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_A = CLBLL_L_X2Y174_SLICE_X1Y174_AO6;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_B = CLBLL_L_X2Y174_SLICE_X1Y174_BO6;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_C = CLBLL_L_X2Y174_SLICE_X1Y174_CO6;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_D = CLBLL_L_X2Y174_SLICE_X1Y174_DO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A = CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B = CLBLL_L_X2Y175_SLICE_X0Y175_BO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C = CLBLL_L_X2Y175_SLICE_X0Y175_CO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D = CLBLL_L_X2Y175_SLICE_X0Y175_DO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A = CLBLL_L_X2Y175_SLICE_X1Y175_AO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B = CLBLL_L_X2Y175_SLICE_X1Y175_BO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C = CLBLL_L_X2Y175_SLICE_X1Y175_CO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D = CLBLL_L_X2Y175_SLICE_X1Y175_DO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A = CLBLL_L_X102Y125_SLICE_X160Y125_AO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B = CLBLL_L_X102Y125_SLICE_X160Y125_BO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C = CLBLL_L_X102Y125_SLICE_X160Y125_CO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D = CLBLL_L_X102Y125_SLICE_X160Y125_DO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A = CLBLL_L_X102Y125_SLICE_X161Y125_AO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B = CLBLL_L_X102Y125_SLICE_X161Y125_BO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C = CLBLL_L_X102Y125_SLICE_X161Y125_CO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D = CLBLL_L_X102Y125_SLICE_X161Y125_DO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_A = CLBLL_R_X81Y111_SLICE_X126Y111_AO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_B = CLBLL_R_X81Y111_SLICE_X126Y111_BO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_C = CLBLL_R_X81Y111_SLICE_X126Y111_CO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_D = CLBLL_R_X81Y111_SLICE_X126Y111_DO6;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_A = CLBLL_R_X81Y111_SLICE_X127Y111_AO6;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_B = CLBLL_R_X81Y111_SLICE_X127Y111_BO6;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_C = CLBLL_R_X81Y111_SLICE_X127Y111_CO6;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_D = CLBLL_R_X81Y111_SLICE_X127Y111_DO6;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_A = CLBLL_R_X81Y122_SLICE_X126Y122_AO6;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_B = CLBLL_R_X81Y122_SLICE_X126Y122_BO6;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_C = CLBLL_R_X81Y122_SLICE_X126Y122_CO6;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_D = CLBLL_R_X81Y122_SLICE_X126Y122_DO6;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_A = CLBLL_R_X81Y122_SLICE_X127Y122_AO6;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_B = CLBLL_R_X81Y122_SLICE_X127Y122_BO6;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_C = CLBLL_R_X81Y122_SLICE_X127Y122_CO6;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_D = CLBLL_R_X81Y122_SLICE_X127Y122_DO6;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_A = CLBLL_R_X81Y124_SLICE_X126Y124_AO6;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_B = CLBLL_R_X81Y124_SLICE_X126Y124_BO6;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_C = CLBLL_R_X81Y124_SLICE_X126Y124_CO6;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_D = CLBLL_R_X81Y124_SLICE_X126Y124_DO6;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_A = CLBLL_R_X81Y124_SLICE_X127Y124_AO6;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_B = CLBLL_R_X81Y124_SLICE_X127Y124_BO6;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_C = CLBLL_R_X81Y124_SLICE_X127Y124_CO6;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_D = CLBLL_R_X81Y124_SLICE_X127Y124_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_AMUX = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_AMUX = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_BMUX = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_CMUX = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_AMUX = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_CMUX = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_DMUX = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_AMUX = CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_A = CLBLM_L_X30Y111_SLICE_X44Y111_AO6;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_B = CLBLM_L_X30Y111_SLICE_X44Y111_BO6;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_C = CLBLM_L_X30Y111_SLICE_X44Y111_CO6;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_D = CLBLM_L_X30Y111_SLICE_X44Y111_DO6;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_A = CLBLM_L_X30Y111_SLICE_X45Y111_AO6;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_B = CLBLM_L_X30Y111_SLICE_X45Y111_BO6;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_C = CLBLM_L_X30Y111_SLICE_X45Y111_CO6;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_D = CLBLM_L_X30Y111_SLICE_X45Y111_DO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_A = CLBLM_L_X46Y121_SLICE_X70Y121_AO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_B = CLBLM_L_X46Y121_SLICE_X70Y121_BO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_C = CLBLM_L_X46Y121_SLICE_X70Y121_CO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_D = CLBLM_L_X46Y121_SLICE_X70Y121_DO6;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_A = CLBLM_L_X46Y121_SLICE_X71Y121_AO6;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_B = CLBLM_L_X46Y121_SLICE_X71Y121_BO6;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_C = CLBLM_L_X46Y121_SLICE_X71Y121_CO6;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_D = CLBLM_L_X46Y121_SLICE_X71Y121_DO6;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_A = CLBLM_L_X46Y142_SLICE_X70Y142_AO6;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_B = CLBLM_L_X46Y142_SLICE_X70Y142_BO6;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_C = CLBLM_L_X46Y142_SLICE_X70Y142_CO6;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_D = CLBLM_L_X46Y142_SLICE_X70Y142_DO6;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_A = CLBLM_L_X46Y142_SLICE_X71Y142_AO6;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_B = CLBLM_L_X46Y142_SLICE_X71Y142_BO6;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_C = CLBLM_L_X46Y142_SLICE_X71Y142_CO6;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_D = CLBLM_L_X46Y142_SLICE_X71Y142_DO6;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_A = CLBLM_L_X50Y119_SLICE_X76Y119_AO6;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_B = CLBLM_L_X50Y119_SLICE_X76Y119_BO6;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_C = CLBLM_L_X50Y119_SLICE_X76Y119_CO6;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_D = CLBLM_L_X50Y119_SLICE_X76Y119_DO6;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_AMUX = CLBLM_L_X50Y119_SLICE_X76Y119_AO5;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_A = CLBLM_L_X50Y119_SLICE_X77Y119_AO6;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_B = CLBLM_L_X50Y119_SLICE_X77Y119_BO6;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_C = CLBLM_L_X50Y119_SLICE_X77Y119_CO6;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_D = CLBLM_L_X50Y119_SLICE_X77Y119_DO6;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D = CLBLM_L_X78Y119_SLICE_X120Y119_DO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A = CLBLM_L_X78Y119_SLICE_X121Y119_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B = CLBLM_L_X78Y119_SLICE_X121Y119_BO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C = CLBLM_L_X78Y119_SLICE_X121Y119_CO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D = CLBLM_L_X78Y119_SLICE_X121Y119_DO6;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_A = CLBLM_L_X78Y125_SLICE_X120Y125_AO6;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_B = CLBLM_L_X78Y125_SLICE_X120Y125_BO6;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_C = CLBLM_L_X78Y125_SLICE_X120Y125_CO6;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_D = CLBLM_L_X78Y125_SLICE_X120Y125_DO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_A = CLBLM_L_X78Y125_SLICE_X121Y125_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_B = CLBLM_L_X78Y125_SLICE_X121Y125_BO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_C = CLBLM_L_X78Y125_SLICE_X121Y125_CO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_D = CLBLM_L_X78Y125_SLICE_X121Y125_DO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A = CLBLM_L_X92Y125_SLICE_X144Y125_AO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B = CLBLM_L_X92Y125_SLICE_X144Y125_BO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C = CLBLM_L_X92Y125_SLICE_X144Y125_CO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D = CLBLM_L_X92Y125_SLICE_X144Y125_DO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_AMUX = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_BMUX = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A = CLBLM_L_X92Y125_SLICE_X145Y125_AO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B = CLBLM_L_X92Y125_SLICE_X145Y125_BO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C = CLBLM_L_X92Y125_SLICE_X145Y125_CO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D = CLBLM_L_X92Y125_SLICE_X145Y125_DO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A = CLBLM_L_X94Y122_SLICE_X148Y122_AO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B = CLBLM_L_X94Y122_SLICE_X148Y122_BO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C = CLBLM_L_X94Y122_SLICE_X148Y122_CO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D = CLBLM_L_X94Y122_SLICE_X148Y122_DO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A = CLBLM_L_X94Y122_SLICE_X149Y122_AO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B = CLBLM_L_X94Y122_SLICE_X149Y122_BO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C = CLBLM_L_X94Y122_SLICE_X149Y122_CO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D = CLBLM_L_X94Y122_SLICE_X149Y122_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_AMUX = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_AMUX = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_AMUX = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_DMUX = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_AMUX = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_BMUX = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_CMUX = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_AMUX = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_AMUX = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_AMUX = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_AMUX = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_BMUX = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AMUX = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_BMUX = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_AMUX = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B = CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C = CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B = CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C = CLBLM_R_X13Y109_SLICE_X19Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D = CLBLM_R_X13Y109_SLICE_X19Y109_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A = CLBLM_R_X13Y110_SLICE_X18Y110_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B = CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C = CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A = CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D = CLBLM_R_X13Y110_SLICE_X19Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_AMUX = CLBLM_R_X13Y110_SLICE_X19Y110_AO5;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_BMUX = CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A = CLBLM_R_X13Y111_SLICE_X18Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B = CLBLM_R_X13Y111_SLICE_X18Y111_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B = CLBLM_R_X13Y111_SLICE_X19Y111_BO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C = CLBLM_R_X13Y111_SLICE_X19Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D = CLBLM_R_X13Y111_SLICE_X19Y111_DO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_AMUX = CLBLM_R_X13Y111_SLICE_X19Y111_AO5;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A = CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B = CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C = CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D = CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_AMUX = CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B = CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C = CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A = CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B = CLBLM_R_X13Y113_SLICE_X18Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C = CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A = CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D = CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_AMUX = CLBLM_R_X13Y113_SLICE_X19Y113_AO5;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_BMUX = CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_A = CLBLM_R_X15Y99_SLICE_X20Y99_AO6;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_B = CLBLM_R_X15Y99_SLICE_X20Y99_BO6;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_C = CLBLM_R_X15Y99_SLICE_X20Y99_CO6;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_D = CLBLM_R_X15Y99_SLICE_X20Y99_DO6;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_AMUX = CLBLM_R_X15Y99_SLICE_X20Y99_AO5;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_A = CLBLM_R_X15Y99_SLICE_X21Y99_AO6;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_B = CLBLM_R_X15Y99_SLICE_X21Y99_BO6;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_C = CLBLM_R_X15Y99_SLICE_X21Y99_CO6;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_D = CLBLM_R_X15Y99_SLICE_X21Y99_DO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A = CLBLM_R_X15Y101_SLICE_X20Y101_AO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B = CLBLM_R_X15Y101_SLICE_X20Y101_BO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C = CLBLM_R_X15Y101_SLICE_X20Y101_CO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D = CLBLM_R_X15Y101_SLICE_X20Y101_DO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_AMUX = CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A = CLBLM_R_X15Y101_SLICE_X21Y101_AO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B = CLBLM_R_X15Y101_SLICE_X21Y101_BO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C = CLBLM_R_X15Y101_SLICE_X21Y101_CO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D = CLBLM_R_X15Y101_SLICE_X21Y101_DO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A = CLBLM_R_X15Y109_SLICE_X20Y109_AO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B = CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C = CLBLM_R_X15Y109_SLICE_X20Y109_CO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D = CLBLM_R_X15Y109_SLICE_X20Y109_DO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_AMUX = CLBLM_R_X15Y109_SLICE_X20Y109_AO5;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A = CLBLM_R_X15Y109_SLICE_X21Y109_AO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B = CLBLM_R_X15Y109_SLICE_X21Y109_BO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C = CLBLM_R_X15Y109_SLICE_X21Y109_CO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D = CLBLM_R_X15Y109_SLICE_X21Y109_DO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A = CLBLM_R_X15Y110_SLICE_X20Y110_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B = CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C = CLBLM_R_X15Y110_SLICE_X20Y110_CO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D = CLBLM_R_X15Y110_SLICE_X20Y110_DO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_AMUX = CLBLM_R_X15Y110_SLICE_X20Y110_AO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A = CLBLM_R_X15Y110_SLICE_X21Y110_AO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B = CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C = CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D = CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_AMUX = CLBLM_R_X15Y110_SLICE_X21Y110_AO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_BMUX = CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A = CLBLM_R_X15Y111_SLICE_X20Y111_AO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C = CLBLM_R_X15Y111_SLICE_X20Y111_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D = CLBLM_R_X15Y111_SLICE_X20Y111_DO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A = CLBLM_R_X15Y111_SLICE_X21Y111_AO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B = CLBLM_R_X15Y111_SLICE_X21Y111_BO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C = CLBLM_R_X15Y111_SLICE_X21Y111_CO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D = CLBLM_R_X15Y111_SLICE_X21Y111_DO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_AMUX = CLBLM_R_X15Y111_SLICE_X21Y111_AO5;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A = CLBLM_R_X15Y113_SLICE_X20Y113_AO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B = CLBLM_R_X15Y113_SLICE_X20Y113_BO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D = CLBLM_R_X15Y113_SLICE_X20Y113_DO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_AMUX = CLBLM_R_X15Y113_SLICE_X20Y113_AO5;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_BMUX = CLBLM_R_X15Y113_SLICE_X20Y113_BO5;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B = CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C = CLBLM_R_X15Y113_SLICE_X21Y113_CO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D = CLBLM_R_X15Y113_SLICE_X21Y113_DO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_AMUX = CLBLM_R_X15Y113_SLICE_X21Y113_AO5;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_BMUX = CLBLM_R_X15Y113_SLICE_X21Y113_BO5;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A = CLBLM_R_X15Y114_SLICE_X20Y114_AO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B = CLBLM_R_X15Y114_SLICE_X20Y114_BO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C = CLBLM_R_X15Y114_SLICE_X20Y114_CO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_AMUX = CLBLM_R_X15Y114_SLICE_X20Y114_AO5;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_BMUX = CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A = CLBLM_R_X15Y114_SLICE_X21Y114_AO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B = CLBLM_R_X15Y114_SLICE_X21Y114_BO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C = CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D = CLBLM_R_X15Y114_SLICE_X21Y114_DO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B = CLBLM_R_X15Y123_SLICE_X20Y123_BO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C = CLBLM_R_X15Y123_SLICE_X20Y123_CO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D = CLBLM_R_X15Y123_SLICE_X20Y123_DO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A = CLBLM_R_X15Y123_SLICE_X21Y123_AO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B = CLBLM_R_X15Y123_SLICE_X21Y123_BO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C = CLBLM_R_X15Y123_SLICE_X21Y123_CO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D = CLBLM_R_X15Y123_SLICE_X21Y123_DO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_A = CLBLM_R_X37Y111_SLICE_X56Y111_AO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_B = CLBLM_R_X37Y111_SLICE_X56Y111_BO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_C = CLBLM_R_X37Y111_SLICE_X56Y111_CO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_D = CLBLM_R_X37Y111_SLICE_X56Y111_DO6;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_A = CLBLM_R_X37Y111_SLICE_X57Y111_AO6;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_B = CLBLM_R_X37Y111_SLICE_X57Y111_BO6;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_C = CLBLM_R_X37Y111_SLICE_X57Y111_CO6;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_D = CLBLM_R_X37Y111_SLICE_X57Y111_DO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A = CLBLM_R_X93Y116_SLICE_X146Y116_AO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B = CLBLM_R_X93Y116_SLICE_X146Y116_BO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C = CLBLM_R_X93Y116_SLICE_X146Y116_CO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D = CLBLM_R_X93Y116_SLICE_X146Y116_DO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A = CLBLM_R_X93Y116_SLICE_X147Y116_AO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B = CLBLM_R_X93Y116_SLICE_X147Y116_BO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C = CLBLM_R_X93Y116_SLICE_X147Y116_CO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D = CLBLM_R_X93Y116_SLICE_X147Y116_DO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A = CLBLM_R_X93Y122_SLICE_X146Y122_AO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B = CLBLM_R_X93Y122_SLICE_X146Y122_BO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C = CLBLM_R_X93Y122_SLICE_X146Y122_CO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D = CLBLM_R_X93Y122_SLICE_X146Y122_DO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A = CLBLM_R_X93Y122_SLICE_X147Y122_AO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B = CLBLM_R_X93Y122_SLICE_X147Y122_BO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C = CLBLM_R_X93Y122_SLICE_X147Y122_CO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D = CLBLM_R_X93Y122_SLICE_X147Y122_DO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A = CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B = CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C = CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D = CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_AMUX = CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A = CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B = CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C = CLBLM_R_X101Y123_SLICE_X159Y123_CO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D = CLBLM_R_X101Y123_SLICE_X159Y123_DO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A = CLBLM_R_X101Y124_SLICE_X158Y124_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B = CLBLM_R_X101Y124_SLICE_X158Y124_BO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C = CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D = CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A = CLBLM_R_X101Y124_SLICE_X159Y124_AO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B = CLBLM_R_X101Y124_SLICE_X159Y124_BO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C = CLBLM_R_X101Y124_SLICE_X159Y124_CO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D = CLBLM_R_X101Y124_SLICE_X159Y124_DO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A = CLBLM_R_X103Y97_SLICE_X162Y97_AO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B = CLBLM_R_X103Y97_SLICE_X162Y97_BO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C = CLBLM_R_X103Y97_SLICE_X162Y97_CO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D = CLBLM_R_X103Y97_SLICE_X162Y97_DO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A = CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B = CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C = CLBLM_R_X103Y97_SLICE_X163Y97_CO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D = CLBLM_R_X103Y97_SLICE_X163Y97_DO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_A = CLBLM_R_X103Y103_SLICE_X162Y103_AO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_B = CLBLM_R_X103Y103_SLICE_X162Y103_BO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_C = CLBLM_R_X103Y103_SLICE_X162Y103_CO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_D = CLBLM_R_X103Y103_SLICE_X162Y103_DO6;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_A = CLBLM_R_X103Y103_SLICE_X163Y103_AO6;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_B = CLBLM_R_X103Y103_SLICE_X163Y103_BO6;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_C = CLBLM_R_X103Y103_SLICE_X163Y103_CO6;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_D = CLBLM_R_X103Y103_SLICE_X163Y103_DO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A = CLBLM_R_X103Y107_SLICE_X162Y107_AO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B = CLBLM_R_X103Y107_SLICE_X162Y107_BO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C = CLBLM_R_X103Y107_SLICE_X162Y107_CO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D = CLBLM_R_X103Y107_SLICE_X162Y107_DO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A = CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B = CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C = CLBLM_R_X103Y107_SLICE_X163Y107_CO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D = CLBLM_R_X103Y107_SLICE_X163Y107_DO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_AMUX = CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A = CLBLM_R_X103Y108_SLICE_X162Y108_AO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B = CLBLM_R_X103Y108_SLICE_X162Y108_BO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C = CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D = CLBLM_R_X103Y108_SLICE_X162Y108_DO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B = CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C = CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D = CLBLM_R_X103Y108_SLICE_X163Y108_DO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_AMUX = CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A = CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B = CLBLM_R_X103Y122_SLICE_X162Y122_BO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C = CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D = CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B = CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C = CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A = CLBLM_R_X103Y125_SLICE_X162Y125_AO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B = CLBLM_R_X103Y125_SLICE_X162Y125_BO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C = CLBLM_R_X103Y125_SLICE_X162Y125_CO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D = CLBLM_R_X103Y125_SLICE_X162Y125_DO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A = CLBLM_R_X103Y125_SLICE_X163Y125_AO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B = CLBLM_R_X103Y125_SLICE_X163Y125_BO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C = CLBLM_R_X103Y125_SLICE_X163Y125_CO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D = CLBLM_R_X103Y125_SLICE_X163Y125_DO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_AMUX = CLBLM_R_X103Y125_SLICE_X163Y125_AO5;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A = CLBLM_R_X103Y147_SLICE_X162Y147_AO6;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B = CLBLM_R_X103Y147_SLICE_X162Y147_BO6;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C = CLBLM_R_X103Y147_SLICE_X162Y147_CO6;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D = CLBLM_R_X103Y147_SLICE_X162Y147_DO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A = CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B = CLBLM_R_X103Y147_SLICE_X163Y147_BO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C = CLBLM_R_X103Y147_SLICE_X163Y147_CO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D = CLBLM_R_X103Y147_SLICE_X163Y147_DO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_AMUX = CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A = CLBLM_R_X103Y185_SLICE_X162Y185_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B = CLBLM_R_X103Y185_SLICE_X162Y185_BO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C = CLBLM_R_X103Y185_SLICE_X162Y185_CO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D = CLBLM_R_X103Y185_SLICE_X162Y185_DO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A = CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B = CLBLM_R_X103Y185_SLICE_X163Y185_BO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C = CLBLM_R_X103Y185_SLICE_X163Y185_CO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D = CLBLM_R_X103Y185_SLICE_X163Y185_DO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_O = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_O = LIOB33_X0Y83_IOB_X0Y84_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_O = LIOB33_X0Y83_IOB_X0Y83_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y86_O = LIOB33_X0Y85_IOB_X0Y86_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y90_O = LIOB33_X0Y89_IOB_X0Y90_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y89_O = LIOB33_X0Y89_IOB_X0Y89_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y92_O = LIOB33_X0Y91_IOB_X0Y92_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y91_O = LIOB33_X0Y91_IOB_X0Y91_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y96_O = LIOB33_X0Y95_IOB_X0Y96_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y95_O = LIOB33_X0Y95_IOB_X0Y95_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y98_O = LIOB33_X0Y97_IOB_X0Y98_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y97_O = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_O = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_O = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_O = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_O = LIOB33_X0Y139_IOB_X0Y140_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_O = LIOB33_X0Y139_IOB_X0Y139_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_O = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_O = LIOB33_X0Y141_IOB_X0Y141_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_O = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_O = LIOB33_X0Y145_IOB_X0Y145_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_O = LIOB33_X0Y147_IOB_X0Y147_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_O = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_O = LIOB33_X0Y151_IOB_X0Y151_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_O = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_O = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_O = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_O = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_O = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_O = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_O = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_O = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_O = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_O = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_O = LIOB33_X0Y171_IOB_X0Y171_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_O = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_O = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_O = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_O = LIOB33_X0Y175_IOB_X0Y175_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_O = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = 1'b0;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = CLBLL_L_X2Y101_SLICE_X0Y101_BO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y99_ILOGIC_X0Y99_O = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_O = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_OQ = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_O = LIOB33_X0Y93_IOB_X0Y94_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_O = LIOB33_X0Y93_IOB_X0Y93_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O = LIOB33_X0Y119_IOB_X0Y119_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O = LIOB33_X0Y131_IOB_X0Y131_I;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O = LIOB33_X0Y143_IOB_X0Y143_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_O = LIOB33_X0Y87_IOB_X0Y88_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_O = LIOB33_X0Y87_IOB_X0Y87_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_O = LIOB33_X0Y137_IOB_X0Y138_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O = LIOB33_X0Y163_IOB_X0Y164_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O = LIOB33_X0Y163_IOB_X0Y163_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_OQ = CLBLM_R_X15Y99_SLICE_X20Y99_AO6;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_OQ = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_OQ = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_OQ = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_OQ = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_OQ = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_OQ = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_OQ = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_OQ = CLBLL_R_X81Y122_SLICE_X126Y122_BO6;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_OQ = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_OQ = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_OQ = CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_OQ = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_OQ = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_OQ = CLBLM_L_X92Y125_SLICE_X144Y125_BO6;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_OQ = CLBLM_L_X92Y125_SLICE_X144Y125_AO6;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_OQ = CLBLL_R_X81Y111_SLICE_X126Y111_AO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_OQ = CLBLM_R_X37Y111_SLICE_X56Y111_BO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_OQ = CLBLM_R_X37Y111_SLICE_X56Y111_CO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_OQ = CLBLM_L_X30Y111_SLICE_X44Y111_AO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_OQ = CLBLL_R_X81Y111_SLICE_X126Y111_BO6;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_TQ = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_OQ = CLBLM_R_X37Y111_SLICE_X56Y111_DO6;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_OQ = CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_OQ = CLBLM_L_X30Y111_SLICE_X44Y111_BO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_OQ = CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_OQ = CLBLM_R_X103Y103_SLICE_X163Y103_AO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_OQ = CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_OQ = CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_OQ = CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_OQ = CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_OQ = CLBLM_R_X15Y113_SLICE_X21Y113_CO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_OQ = CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_OQ = CLBLM_R_X15Y113_SLICE_X20Y113_DO6;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_OQ = CLBLM_R_X15Y114_SLICE_X20Y114_CO6;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_OQ = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_OQ = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_OQ = CLBLL_L_X102Y125_SLICE_X161Y125_AO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLM_R_X37Y111_SLICE_X56Y111_AO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLM_R_X101Y124_SLICE_X158Y124_AO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLL_L_X102Y125_SLICE_X161Y125_BO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLM_R_X93Y122_SLICE_X147Y122_CO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_R_X101Y124_SLICE_X158Y124_BO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = CLBLM_L_X94Y122_SLICE_X148Y122_AO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLM_L_X78Y119_SLICE_X121Y119_CO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLM_L_X94Y122_SLICE_X148Y122_BO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = CLBLM_L_X78Y119_SLICE_X121Y119_DO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLM_R_X103Y125_SLICE_X162Y125_BO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = CLBLM_L_X78Y125_SLICE_X121Y125_BO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLM_L_X78Y125_SLICE_X121Y125_AO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLM_L_X78Y125_SLICE_X121Y125_DO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLM_L_X78Y125_SLICE_X121Y125_CO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_X105Y151_ILOGIC_X1Y152_O = RIOB33_X105Y151_IOB_X1Y152_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y151_O = RIOB33_X105Y151_IOB_X1Y151_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y154_O = RIOB33_X105Y153_IOB_X1Y154_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y153_O = RIOB33_X105Y153_IOB_X1Y153_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y156_O = RIOB33_X105Y155_IOB_X1Y156_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y155_O = RIOB33_X105Y155_IOB_X1Y155_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y160_O = RIOB33_X105Y159_IOB_X1Y160_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y159_O = RIOB33_X105Y159_IOB_X1Y159_I;
  assign RIOI3_X105Y161_ILOGIC_X1Y161_O = RIOB33_X105Y161_IOB_X1Y161_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y166_O = RIOB33_X105Y165_IOB_X1Y166_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y165_O = RIOB33_X105Y165_IOB_X1Y165_I;
  assign RIOI3_X105Y167_ILOGIC_X1Y168_O = RIOB33_X105Y167_IOB_X1Y168_I;
  assign RIOI3_X105Y167_ILOGIC_X1Y167_O = RIOB33_X105Y167_IOB_X1Y167_I;
  assign RIOI3_X105Y171_ILOGIC_X1Y172_O = RIOB33_X105Y171_IOB_X1Y172_I;
  assign RIOI3_X105Y171_ILOGIC_X1Y171_O = RIOB33_X105Y171_IOB_X1Y171_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = LIOB33_X0Y133_IOB_X0Y133_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = LIOB33_X0Y137_IOB_X0Y138_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = LIOB33_X0Y103_IOB_X0Y104_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = LIOB33_X0Y133_IOB_X0Y134_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLL_L_X2Y174_SLICE_X0Y174_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLL_L_X2Y174_SLICE_X0Y174_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLL_L_X2Y174_SLICE_X0Y174_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ = CLBLM_R_X15Y99_SLICE_X20Y99_AO6;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ = CLBLM_L_X78Y119_SLICE_X121Y119_BO6;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_SING_X105Y150_ILOGIC_X1Y150_O = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLL_L_X2Y174_SLICE_X0Y174_BO5;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ = CLBLL_R_X81Y122_SLICE_X126Y122_AO6;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ = CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ = CLBLM_R_X15Y110_SLICE_X20Y110_CO6;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ = CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ = CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ = CLBLM_R_X15Y113_SLICE_X21Y113_DO6;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLM_L_X78Y119_SLICE_X121Y119_AO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLM_R_X93Y122_SLICE_X147Y122_AO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_O = RIOB33_X105Y157_IOB_X1Y158_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_O = RIOB33_X105Y157_IOB_X1Y157_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_O = RIOB33_X105Y169_IOB_X1Y170_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_O = RIOB33_X105Y169_IOB_X1Y169_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ = CLBLM_R_X15Y110_SLICE_X20Y110_DO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ = CLBLM_R_X103Y103_SLICE_X163Y103_BO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = CLBLM_R_X103Y125_SLICE_X162Y125_AO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_O = RIOB33_X105Y163_IOB_X1Y163_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y176_O = LIOB33_X0Y137_IOB_X0Y138_I;
  assign RIOB33_X105Y175_IOB_X1Y175_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_D = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = RIOB33_X105Y169_IOB_X1Y170_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLM_L_X94Y122_SLICE_X148Y122_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_D1 = CLBLL_R_X81Y111_SLICE_X126Y111_BO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_T1 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = CLBLM_L_X78Y119_SLICE_X121Y119_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_D1 = CLBLM_R_X37Y111_SLICE_X56Y111_DO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = CLBLM_R_X103Y125_SLICE_X162Y125_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign RIOB33_X105Y57_IOB_X1Y58_O = CLBLL_R_X81Y122_SLICE_X126Y122_AO6;
  assign RIOB33_X105Y57_IOB_X1Y57_O = CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C3 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C4 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C5 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A3 = 1'b1;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_D = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_D = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOB33_X105Y177_IOB_X1Y177_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A4 = 1'b1;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLL_L_X2Y174_SLICE_X0Y174_BO5;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D2 = 1'b1;
  assign LIOI3_X0Y95_ILOGIC_X0Y96_D = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D3 = 1'b1;
  assign LIOI3_X0Y95_ILOGIC_X0Y95_D = LIOB33_X0Y95_IOB_X0Y95_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign RIOI3_X105Y171_ILOGIC_X1Y172_D = RIOB33_X105Y171_IOB_X1Y172_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D4 = 1'b1;
  assign RIOI3_X105Y171_ILOGIC_X1Y171_D = RIOB33_X105Y171_IOB_X1Y171_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D5 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A5 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A1 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A3 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A4 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A5 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A2 = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A4 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B1 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B2 = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B4 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B6 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D4 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D5 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A5 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A1 = CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A2 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A5 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_A1 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_A2 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_A3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_A4 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_A5 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_B1 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_B2 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_B3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_B4 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_B5 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_B6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_C1 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_C2 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_C3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_C4 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_C5 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_D1 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_D2 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_D3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_D4 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_L_X50Y119_SLICE_X77Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_A1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_A2 = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_A3 = CLBLM_R_X15Y113_SLICE_X21Y113_DO6;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_A4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_A6 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_B1 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_B2 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_B3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_B4 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_B5 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_B6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_C1 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_C2 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_C3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_C4 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_C5 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B1 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_D1 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_D2 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_D3 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_D4 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_D5 = 1'b1;
  assign CLBLM_L_X50Y119_SLICE_X76Y119_D6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B3 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D3 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D4 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D5 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B4 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B5 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A6 = 1'b1;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_B2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B1 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B2 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B4 = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B6 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A1 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A2 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A3 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A4 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A5 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C2 = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B1 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B2 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B4 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B5 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C1 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C2 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D1 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D2 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D3 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D4 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D5 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A1 = CLBLM_R_X15Y113_SLICE_X20Y113_BO5;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A3 = CLBLL_R_X81Y124_SLICE_X126Y124_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A5 = CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A6 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A1 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A2 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A4 = CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A5 = LIOB33_X0Y89_IOB_X0Y90_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A6 = CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B1 = CLBLM_R_X15Y113_SLICE_X20Y113_BO5;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B2 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B3 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B4 = CLBLL_R_X81Y122_SLICE_X126Y122_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B1 = LIOB33_X0Y87_IOB_X0Y87_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B2 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B3 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B4 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B5 = LIOB33_X0Y91_IOB_X0Y92_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B6 = CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C2 = CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C3 = CLBLM_R_X15Y113_SLICE_X20Y113_BO5;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C4 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C5 = CLBLM_R_X13Y110_SLICE_X19Y110_AO5;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D2 = CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D3 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D4 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D5 = CLBLM_R_X15Y113_SLICE_X20Y113_BO5;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D2 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D3 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D5 = LIOB33_X0Y87_IOB_X0Y87_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D6 = 1'b1;
  assign RIOB33_X105Y61_IOB_X1Y61_O = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign RIOB33_X105Y61_IOB_X1Y62_O = CLBLL_R_X81Y122_SLICE_X126Y122_BO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C2 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C3 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C4 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLM_R_X103Y125_SLICE_X162Y125_BO6;
  assign RIOB33_X105Y181_IOB_X1Y182_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_D1 = CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C5 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_D1 = CLBLM_R_X15Y99_SLICE_X20Y99_AO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_D1 = CLBLM_L_X30Y111_SLICE_X44Y111_BO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C6 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_D1 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1 = CLBLL_R_X81Y122_SLICE_X126Y122_AO6;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1 = CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B1 = LIOB33_X0Y93_IOB_X0Y94_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B2 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B3 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C1 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C5 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C6 = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_D = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D6 = 1'b1;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_D = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A6 = 1'b1;
  assign LIOI3_X0Y97_ILOGIC_X0Y98_D = LIOB33_X0Y97_IOB_X0Y98_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y97_D = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B6 = 1'b1;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOB33_X105Y63_IOB_X1Y63_O = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign RIOB33_X105Y63_IOB_X1Y64_O = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C3 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C4 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C5 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C6 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_D = RIOB33_X105Y163_IOB_X1Y163_I;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_A1 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_A2 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_A3 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_A4 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_A5 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_A6 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_B1 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_B2 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_B3 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_B4 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_B5 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_B6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D1 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y183_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOB33_X105Y183_IOB_X1Y184_O = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_C1 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_C2 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_C3 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_C4 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_C5 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_C6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_D = LIOB33_X0Y93_IOB_X0Y94_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D4 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_D1 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_D2 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_D3 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_D4 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_D5 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X45Y111_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_D = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_A1 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_A2 = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_A3 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_A4 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_A5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_A6 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_B1 = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_B2 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_B3 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_B4 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_B5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_B6 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_C1 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_C2 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_C3 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_C4 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_C5 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_C6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A1 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_D1 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_D2 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_D3 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_D4 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_D5 = 1'b1;
  assign CLBLM_L_X30Y111_SLICE_X44Y111_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A1 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A4 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A5 = LIOB33_X0Y91_IOB_X0Y92_I;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C1 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B1 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B2 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B4 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C1 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C2 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C4 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C5 = 1'b1;
  assign RIOB33_X105Y65_IOB_X1Y65_O = CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  assign RIOB33_X105Y65_IOB_X1Y66_O = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_C3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D1 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D2 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D4 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_C4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_C5 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A2 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A3 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A1 = CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A2 = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A4 = CLBLM_R_X13Y111_SLICE_X18Y111_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A5 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A6 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A4 = CLBLM_R_X93Y122_SLICE_X147Y122_BO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A5 = CLBLL_R_X81Y124_SLICE_X126Y124_AO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B1 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B5 = LIOB33_X0Y91_IOB_X0Y92_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B6 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B2 = RIOB33_X105Y151_IOB_X1Y151_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B3 = CLBLM_R_X15Y111_SLICE_X21Y111_BO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B4 = RIOB33_X105Y151_IOB_X1Y152_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B6 = CLBLM_R_X15Y113_SLICE_X20Y113_AO5;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_A1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_A2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_A3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C6 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_A4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_A5 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_A6 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C2 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_B1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_B2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_B3 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_B4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_B5 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_B6 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D1 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_C1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_C2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_C3 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_C4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_C5 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_C6 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D6 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D4 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A5 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A6 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D5 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_D1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_D2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_D3 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_D4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_D5 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X71Y142_D6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B1 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B3 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B4 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B5 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B6 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_A1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_A2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_A3 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_A4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_A5 = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_A6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C3 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C4 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C6 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_B1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_B2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_B3 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_B4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_B5 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_B6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D1 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D3 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_C1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_C2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_C3 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_C4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_C5 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_C6 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_D1 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_D2 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_D3 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_D4 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_D5 = 1'b1;
  assign CLBLM_L_X46Y142_SLICE_X70Y142_D6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_A5 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_A6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLL_L_X2Y174_SLICE_X0Y174_AO5;
  assign RIOI3_X105Y165_ILOGIC_X1Y165_D = RIOB33_X105Y165_IOB_X1Y165_I;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_B3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_B4 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_A3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_A4 = RIOB33_X105Y155_IOB_X1Y155_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_A5 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_A6 = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_B5 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_B6 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_B1 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_B3 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_B4 = RIOB33_X105Y155_IOB_X1Y155_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_B5 = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_B6 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_C1 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_C2 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_C3 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_C4 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_C5 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_C6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_D1 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_D2 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_D3 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_D4 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_D5 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X126Y122_D6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_C1 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_C2 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_C3 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = CLBLM_L_X78Y125_SLICE_X121Y125_BO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_C4 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_C5 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_C6 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_D1 = CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_A1 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_A2 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_A3 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_A4 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_A5 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_A6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A2 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A3 = CLBLM_R_X15Y111_SLICE_X21Y111_AO5;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_B1 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_B2 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_B3 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_B4 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_B5 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_B6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A4 = CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A5 = CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_C1 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_C2 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_C3 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_C4 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_C5 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_C6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B3 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B4 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B6 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_D1 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_D2 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_D3 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_D4 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_D5 = 1'b1;
  assign CLBLL_R_X81Y122_SLICE_X127Y122_D6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D1 = RIOB33_X105Y163_IOB_X1Y163_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D6 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D3 = CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_D1 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLM_R_X37Y111_SLICE_X56Y111_AO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_D2 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y128_O = CLBLL_L_X102Y125_SLICE_X161Y125_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A1 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A2 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A3 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_D3 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_D4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B3 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B4 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A6 = CLBLM_R_X15Y113_SLICE_X20Y113_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_D5 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_D6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C1 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C3 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C5 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C6 = CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D1 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D2 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D3 = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D4 = CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D6 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C2 = 1'b1;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_D = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_D = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_D = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_D = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D = LIOB33_X0Y143_IOB_X0Y143_I;
  assign RIOB33_X105Y69_IOB_X1Y70_O = CLBLM_R_X15Y110_SLICE_X20Y110_CO6;
  assign RIOB33_X105Y69_IOB_X1Y69_O = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A1 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A2 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A3 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A4 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A5 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B1 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B2 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B3 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B4 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B5 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B6 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A2 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C1 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C2 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B1 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B4 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D1 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C1 = CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C2 = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C3 = RIOB33_X105Y171_IOB_X1Y171_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C4 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C5 = CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C6 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D3 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D4 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D5 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A1 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A2 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A3 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D1 = CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D2 = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D3 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D4 = CLBLM_R_X13Y113_SLICE_X19Y113_AO5;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D5 = CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D6 = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A5 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B1 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B2 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A2 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A6 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C5 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D1 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D2 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D4 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D5 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D6 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D6 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D1 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_A2 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_A3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_A4 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_A5 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_A6 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_B1 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_B2 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_B3 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_B4 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_B5 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_B6 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_C1 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_C2 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_C3 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_C4 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_C5 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_C6 = 1'b1;
  assign RIOB33_X105Y71_IOB_X1Y71_O = CLBLM_L_X92Y125_SLICE_X144Y125_AO6;
  assign RIOB33_X105Y71_IOB_X1Y72_O = CLBLM_L_X92Y125_SLICE_X144Y125_BO6;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_D1 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_D2 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_D3 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_D4 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_D5 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X126Y124_D6 = 1'b1;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLM_L_X78Y119_SLICE_X121Y119_AO6;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLM_R_X93Y122_SLICE_X147Y122_AO6;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_A1 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_A2 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_A3 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_A4 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_A5 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_A6 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_B1 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_B2 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_B3 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_B4 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_B5 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_B6 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_C1 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_C2 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_C3 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_C4 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_C5 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_C6 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_D1 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_D2 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_D3 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_D4 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_D5 = 1'b1;
  assign CLBLL_R_X81Y124_SLICE_X127Y124_D6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = 1'b0;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C2 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLM_L_X78Y125_SLICE_X121Y125_DO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_D1 = CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLM_L_X78Y125_SLICE_X121Y125_CO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A1 = RIOB33_X105Y167_IOB_X1Y167_I;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A2 = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_D1 = CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A4 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_D1 = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A5 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_T1 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1 = CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B1 = CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1 = CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B3 = CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B4 = CLBLM_R_X15Y99_SLICE_X20Y99_AO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B5 = CLBLM_R_X15Y110_SLICE_X21Y110_AO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B6 = RIOB33_X105Y167_IOB_X1Y167_I;
  assign RIOB33_X105Y73_IOB_X1Y74_O = CLBLL_R_X81Y111_SLICE_X126Y111_AO6;
  assign RIOB33_X105Y73_IOB_X1Y73_O = CLBLM_R_X37Y111_SLICE_X56Y111_BO6;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_D = LIOB33_X0Y165_IOB_X0Y166_I;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLM_R_X93Y122_SLICE_X147Y122_CO6;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_R_X101Y124_SLICE_X158Y124_BO6;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_D = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_D = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_D = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_A1 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_A2 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_A3 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_A4 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_A5 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_A6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_B1 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_B2 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_B3 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_B4 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_B5 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_D = LIOB33_X0Y87_IOB_X0Y88_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_D = LIOB33_X0Y87_IOB_X0Y87_I;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_C1 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_C2 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_C3 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_C4 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_C5 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_D1 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_D2 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_D3 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_D4 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_D5 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X21Y99_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B1 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_A1 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_A2 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_A3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_A4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_A5 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_A6 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_B1 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_B2 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_B3 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_B4 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_B5 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_B6 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_C1 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_C2 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_C3 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_C4 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_C5 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_C6 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_D1 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_D2 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_D3 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_D4 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_D5 = 1'b1;
  assign CLBLM_R_X15Y99_SLICE_X20Y99_D6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A2 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A3 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C6 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D6 = 1'b1;
  assign LIOI3_X0Y91_ILOGIC_X0Y92_D = LIOB33_X0Y91_IOB_X0Y92_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D6 = 1'b1;
  assign RIOB33_X105Y75_IOB_X1Y75_O = CLBLM_L_X30Y111_SLICE_X44Y111_AO6;
  assign RIOB33_X105Y75_IOB_X1Y76_O = CLBLM_R_X37Y111_SLICE_X56Y111_CO6;
  assign RIOB33_X105Y135_IOB_X1Y136_O = CLBLM_L_X94Y122_SLICE_X148Y122_AO6;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLM_L_X78Y119_SLICE_X121Y119_CO6;
  assign LIOI3_X0Y91_ILOGIC_X0Y91_D = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A1 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A3 = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A4 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A5 = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A6 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  assign RIOB33_X105Y195_IOB_X1Y195_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C6 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D6 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A6 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B6 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C6 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D6 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_A1 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_A2 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_A3 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_A4 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_A5 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_A6 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_B1 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_B2 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_B3 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_B4 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_B5 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_B6 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_C1 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_C2 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_C3 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_C4 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_C5 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_C6 = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1 = CLBLM_R_X15Y99_SLICE_X20Y99_AO6;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_D1 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_D2 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_D3 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_D4 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_D5 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X71Y121_D6 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_A2 = CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_A3 = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_A4 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_A5 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_A6 = CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_B2 = CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_B3 = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_B4 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_B5 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_B6 = CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_C1 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_C2 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_C3 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_C4 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_C5 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_C6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B1 = CLBLM_R_X15Y113_SLICE_X21Y113_BO5;
  assign RIOB33_X105Y77_IOB_X1Y77_O = CLBLM_R_X37Y111_SLICE_X56Y111_DO6;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_D1 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_D2 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_D3 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_D4 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_D5 = 1'b1;
  assign CLBLM_L_X46Y121_SLICE_X70Y121_D6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = CLBLL_L_X2Y101_SLICE_X0Y101_BO6;
  assign RIOB33_X105Y77_IOB_X1Y78_O = CLBLL_R_X81Y111_SLICE_X126Y111_BO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B5 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign RIOB33_X105Y137_IOB_X1Y138_O = CLBLM_R_X103Y125_SLICE_X162Y125_AO6;
  assign RIOB33_X105Y137_IOB_X1Y137_O = CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C2 = CLBLL_R_X81Y122_SLICE_X126Y122_CO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C5 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_D1 = CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C6 = CLBLM_R_X93Y122_SLICE_X147Y122_BO6;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_D1 = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_T1 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_D1 = CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLL_L_X2Y174_SLICE_X0Y174_AO6;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLL_L_X2Y174_SLICE_X0Y174_AO6;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_D1 = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_A1 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_A2 = LIOB33_X0Y97_IOB_X0Y98_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_A3 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_A4 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_A5 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_A6 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_B2 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_B3 = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_B4 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_B5 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_B6 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_C1 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_C2 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_C3 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_C4 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_C5 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_C6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1 = CLBLM_R_X15Y113_SLICE_X21Y113_DO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_D1 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_D2 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_D3 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_D4 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_D5 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X0Y174_D6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A2 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A3 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A4 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D6 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B2 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B3 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B4 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B6 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C2 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C3 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C4 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C6 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_A1 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_A2 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_A3 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_A4 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_A5 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_A6 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D1 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_B1 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_B2 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D6 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_B3 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_B4 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_B5 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_B6 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D3 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_C1 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_C2 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_C3 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_C4 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A5 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A6 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_C5 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_C6 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A1 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A2 = CLBLM_R_X15Y109_SLICE_X20Y109_AO5;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B2 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B3 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B4 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B6 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_D1 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_D2 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_D3 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C2 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C3 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C4 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C6 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_D6 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D2 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D3 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D4 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D6 = 1'b1;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_D = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_D = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B2 = 1'b1;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y152_D = RIOB33_X105Y151_IOB_X1Y152_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y151_D = RIOB33_X105Y151_IOB_X1Y151_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A2 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A3 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A5 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B2 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B3 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B5 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C2 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C3 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C5 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C6 = 1'b1;
  assign RIOB33_X105Y79_IOB_X1Y79_O = CLBLM_L_X30Y111_SLICE_X44Y111_BO6;
  assign RIOB33_X105Y79_IOB_X1Y80_O = CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A1 = CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A3 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D2 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D3 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D5 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A2 = CLBLM_R_X103Y125_SLICE_X163Y125_AO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A3 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A5 = CLBLL_R_X81Y122_SLICE_X126Y122_CO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A6 = CLBLM_R_X15Y114_SLICE_X20Y114_AO5;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A2 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A3 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A4 = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B2 = CLBLM_R_X103Y125_SLICE_X163Y125_AO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B3 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B4 = CLBLL_R_X81Y124_SLICE_X126Y124_AO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B2 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B3 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B4 = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C2 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D2 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D3 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D5 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D4 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C1 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y192_O = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C3 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y191_O = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A3 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A5 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C5 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_T1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D2 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D4 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A2 = CLBLM_R_X15Y114_SLICE_X20Y114_AO5;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A3 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A4 = CLBLM_R_X103Y125_SLICE_X163Y125_AO5;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A5 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign RIOB33_X105Y81_IOB_X1Y82_O = CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  assign RIOB33_X105Y81_IOB_X1Y81_O = CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B2 = CLBLM_R_X15Y114_SLICE_X20Y114_AO5;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B3 = CLBLM_R_X103Y125_SLICE_X163Y125_AO5;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B6 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLM_R_X103Y125_SLICE_X162Y125_BO6;
  assign RIOB33_X105Y89_IOB_X1Y90_O = CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  assign RIOB33_X105Y89_IOB_X1Y89_O = CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C6 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_D1 = CLBLM_R_X15Y113_SLICE_X21Y113_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOB33_X105Y185_IOB_X1Y186_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOB33_X105Y185_IOB_X1Y185_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = LIOB33_X0Y97_IOB_X0Y97_I;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_D1 = CLBLL_R_X81Y122_SLICE_X126Y122_BO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_T1 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_D1 = CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_D1 = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign RIOB33_X105Y83_IOB_X1Y83_O = CLBLM_R_X103Y103_SLICE_X163Y103_AO6;
  assign RIOB33_X105Y83_IOB_X1Y84_O = CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign RIOB33_X105Y143_IOB_X1Y144_O = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A2 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A3 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A5 = RIOB33_X105Y165_IOB_X1Y165_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A1 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_O = CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_D = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B1 = CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_D = LIOB33_X0Y171_IOB_X0Y171_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_D = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B2 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_D = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B3 = CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B5 = CLBLM_R_X15Y110_SLICE_X20Y110_AO5;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y154_D = RIOB33_X105Y153_IOB_X1Y154_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y153_D = RIOB33_X105Y153_IOB_X1Y153_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C3 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_D = LIOB33_X0Y137_IOB_X0Y138_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A2 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A3 = CLBLL_R_X81Y124_SLICE_X126Y124_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A4 = CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A5 = CLBLM_L_X50Y119_SLICE_X76Y119_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A6 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B1 = CLBLL_R_X81Y122_SLICE_X126Y122_CO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B3 = CLBLM_L_X50Y119_SLICE_X76Y119_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B5 = CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B6 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C1 = CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C2 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C4 = CLBLM_L_X50Y119_SLICE_X76Y119_AO5;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C6 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D1 = CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D4 = CLBLM_L_X50Y119_SLICE_X76Y119_AO5;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D5 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D6 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A2 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A4 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign LIOB33_SING_X0Y200_IOB_X0Y200_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B2 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B4 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C2 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C4 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C6 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D2 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D4 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign RIOB33_X105Y85_IOB_X1Y86_O = CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  assign RIOB33_X105Y85_IOB_X1Y85_O = CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign RIOB33_X105Y145_IOB_X1Y146_O = CLBLM_L_X78Y125_SLICE_X121Y125_BO6;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLM_L_X78Y125_SLICE_X121Y125_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_D1 = CLBLM_L_X92Y125_SLICE_X144Y125_BO6;
  assign LIOB33_X0Y179_IOB_X0Y180_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign RIOB33_X105Y67_IOB_X1Y68_O = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign RIOB33_X105Y67_IOB_X1Y67_O = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D3 = 1'b1;
  assign RIOB33_X105Y87_IOB_X1Y88_O = CLBLM_R_X15Y110_SLICE_X20Y110_DO6;
  assign RIOB33_X105Y87_IOB_X1Y87_O = CLBLM_R_X103Y103_SLICE_X163Y103_BO6;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLM_L_X78Y125_SLICE_X121Y125_DO6;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLM_L_X78Y125_SLICE_X121Y125_CO6;
  assign RIOI3_SING_X105Y150_ILOGIC_X1Y150_D = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOB33_X0Y181_IOB_X0Y181_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_D1 = CLBLM_R_X15Y113_SLICE_X20Y113_DO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_D1 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = 1'b0;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_D1 = CLBLM_R_X15Y114_SLICE_X20Y114_CO6;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_D1 = CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_T1 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLL_L_X2Y174_SLICE_X0Y174_BO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D2 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D4 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLM_R_X101Y124_SLICE_X158Y124_AO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A2 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A4 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A6 = 1'b1;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_D = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B6 = 1'b1;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_D = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_D = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_D = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C6 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_D = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D6 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y156_D = RIOB33_X105Y155_IOB_X1Y156_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y155_D = RIOB33_X105Y155_IOB_X1Y155_I;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D = LIOB33_X0Y163_IOB_X0Y164_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLL_L_X102Y125_SLICE_X161Y125_BO6;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  assign LIOB33_X0Y183_IOB_X0Y183_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOB33_X0Y193_IOB_X0Y194_O = 1'b0;
  assign LIOB33_X0Y193_IOB_X0Y193_O = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_D = LIOB33_X0Y153_IOB_X0Y153_I;
  assign RIOB33_X105Y91_IOB_X1Y92_O = CLBLM_R_X15Y113_SLICE_X21Y113_CO6;
  assign RIOB33_X105Y91_IOB_X1Y91_O = CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A5 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A6 = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_A1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_A3 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_A4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_A5 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_A6 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_B1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_B2 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_B3 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_B4 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_B5 = CLBLL_L_X2Y101_SLICE_X0Y101_AO6;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_B6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_C1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_C2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_C3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_C4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_C5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_C6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B2 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_D1 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_D2 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_D3 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_D4 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_D5 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X0Y101_D6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D6 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_A1 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_A2 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_A3 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_A4 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_A5 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_A6 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_B1 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_B2 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_B3 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_B4 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_B5 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_B6 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_C1 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_C2 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_C3 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_C4 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_C5 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_C6 = 1'b1;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLM_L_X94Y122_SLICE_X148Y122_BO6;
  assign RIOB33_X105Y139_IOB_X1Y139_O = CLBLM_L_X78Y119_SLICE_X121Y119_DO6;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_D1 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_D2 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_D3 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_D4 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_D5 = 1'b1;
  assign CLBLL_L_X2Y101_SLICE_X1Y101_D6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_C6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign RIOI3_X105Y167_ILOGIC_X1Y168_D = RIOB33_X105Y167_IOB_X1Y168_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y167_ILOGIC_X1Y167_D = RIOB33_X105Y167_IOB_X1Y167_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = 1'b1;
  assign RIOB33_X105Y93_IOB_X1Y93_O = CLBLM_R_X15Y113_SLICE_X21Y113_DO6;
  assign RIOB33_X105Y93_IOB_X1Y94_O = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_D1 = CLBLL_L_X102Y125_SLICE_X161Y125_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_D1 = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_T1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_T1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLM_R_X37Y111_SLICE_X56Y111_AO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_T1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_D1 = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A2 = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A4 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A6 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_T1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B2 = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B4 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B6 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLM_R_X93Y122_SLICE_X147Y122_AO6;
  assign LIOB33_X0Y187_IOB_X0Y188_O = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign LIOB33_X0Y187_IOB_X0Y187_O = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D2 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D5 = 1'b1;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_D = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_D = LIOB33_X0Y175_IOB_X0Y175_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_D = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_D = LIOB33_X0Y145_IOB_X0Y145_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D6 = 1'b1;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_D = LIOB33_X0Y83_IOB_X0Y84_I;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1 = CLBLM_R_X15Y110_SLICE_X20Y110_CO6;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_D = LIOB33_X0Y83_IOB_X0Y83_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y160_D = RIOB33_X105Y159_IOB_X1Y160_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y159_D = RIOB33_X105Y159_IOB_X1Y159_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1 = CLBLM_L_X78Y119_SLICE_X121Y119_BO6;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D = LIOB33_X0Y81_IOB_X0Y82_I;
  assign RIOB33_X105Y95_IOB_X1Y96_O = CLBLM_R_X15Y113_SLICE_X20Y113_DO6;
  assign RIOB33_X105Y95_IOB_X1Y95_O = CLBLM_R_X15Y114_SLICE_X20Y114_CO6;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = RIOB33_X105Y169_IOB_X1Y169_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = RIOB33_X105Y167_IOB_X1Y168_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign LIOB33_X0Y189_IOB_X0Y190_O = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign LIOB33_X0Y189_IOB_X0Y189_O = CLBLL_L_X2Y174_SLICE_X0Y174_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A1 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A2 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A3 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A4 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A6 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B2 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B3 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B4 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B6 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C1 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C1 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C2 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C3 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C4 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D1 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D2 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D3 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D4 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C6 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A1 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A2 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A3 = CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A4 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A5 = LIOB33_X0Y93_IOB_X0Y94_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B2 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B3 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B4 = CLBLM_R_X15Y99_SLICE_X20Y99_AO5;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B5 = CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B6 = LIOB33_X0Y93_IOB_X0Y94_I;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C1 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C2 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C3 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C4 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C6 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D1 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D2 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D3 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D4 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A2 = 1'b1;
  assign RIOB33_X105Y97_IOB_X1Y98_O = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign RIOB33_X105Y97_IOB_X1Y97_O = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign RIOI3_X105Y161_ILOGIC_X1Y161_D = RIOB33_X105Y161_IOB_X1Y161_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_A1 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_A2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_A3 = CLBLM_L_X46Y142_SLICE_X70Y142_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_A4 = CLBLL_R_X81Y124_SLICE_X126Y124_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_A5 = CLBLM_L_X46Y121_SLICE_X70Y121_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_A6 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_B3 = CLBLL_R_X81Y122_SLICE_X126Y122_CO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_B4 = CLBLM_L_X46Y121_SLICE_X70Y121_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_B5 = CLBLM_L_X46Y142_SLICE_X70Y142_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_B6 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_B1 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_C1 = CLBLM_L_X46Y142_SLICE_X70Y142_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_C2 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_C3 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_C4 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_C5 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_C6 = CLBLM_L_X46Y121_SLICE_X70Y121_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_D1 = CLBLM_L_X46Y142_SLICE_X70Y142_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_D2 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_D3 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_D4 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_D5 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_L_X78Y125_SLICE_X121Y125_D6 = CLBLM_L_X46Y121_SLICE_X70Y121_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_A1 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_A2 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_A3 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_A4 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_A5 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_A6 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_B1 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_B2 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_B3 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_B4 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_B5 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_B6 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_C1 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_C2 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_C3 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_C4 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_C5 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_C6 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C1 = CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C3 = CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C4 = CLBLM_R_X15Y110_SLICE_X21Y110_AO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C6 = CLBLM_R_X15Y99_SLICE_X20Y99_AO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D1 = CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D2 = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_D1 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_D2 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_D3 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_D4 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_D5 = 1'b1;
  assign CLBLM_L_X78Y125_SLICE_X120Y125_D6 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D3 = CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D4 = CLBLM_R_X15Y111_SLICE_X21Y111_AO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D6 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A4 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A5 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A1 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A2 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A3 = LIOB33_X0Y89_IOB_X0Y90_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A3 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B1 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B2 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B4 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B5 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B6 = CLBLM_R_X15Y111_SLICE_X20Y111_AO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C2 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C3 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C4 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C1 = CLBLM_R_X15Y110_SLICE_X20Y110_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C2 = CLBLM_R_X15Y109_SLICE_X20Y109_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C3 = CLBLM_R_X15Y109_SLICE_X20Y109_AO5;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C4 = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C5 = CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C6 = CLBLM_R_X13Y111_SLICE_X18Y111_AO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A4 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D2 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D3 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D4 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D6 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D1 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D2 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D3 = CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D5 = CLBLM_R_X15Y101_SLICE_X20Y101_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D6 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_T1 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_D1 = CLBLM_L_X92Y125_SLICE_X144Y125_AO6;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLM_R_X101Y124_SLICE_X158Y124_AO6;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_A1 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_A2 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_A3 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_A4 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_A5 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_A6 = 1'b1;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLL_L_X102Y125_SLICE_X161Y125_BO6;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_D = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_B1 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_B2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_B3 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_B4 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_B5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_C1 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_C2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_D1 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_D2 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_D3 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_D4 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_D5 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_A2 = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_A4 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_B1 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_B2 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_B3 = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_B4 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_B5 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_B6 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_C3 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_C5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_C6 = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = RIOB33_X105Y165_IOB_X1Y166_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_D1 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_D2 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_D3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_D4 = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_D5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X37Y111_SLICE_X56Y111_D6 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_A2 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_A3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_A4 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_A5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_A6 = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_B1 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_B2 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_B3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_B4 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_B5 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_B6 = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_C1 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_C2 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_C3 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_C4 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_C5 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_C6 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C1 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C2 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C3 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C4 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C5 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_D1 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D1 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D2 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D3 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D4 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D5 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D6 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_D2 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_D3 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_D4 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_D5 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X126Y111_D6 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A2 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A3 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A5 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A6 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_D1 = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B3 = CLBLM_R_X15Y109_SLICE_X20Y109_AO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B4 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B5 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_D = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_A1 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_A2 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_A3 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_A4 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C4 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C5 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C6 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_A5 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_A6 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C1 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C2 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C3 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_B1 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_B2 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_B3 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_B4 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_B5 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_B6 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D1 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D2 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_C1 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_C2 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_C3 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_C4 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_C5 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_C6 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D4 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D5 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D6 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_D1 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_D2 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_D3 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_D4 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_D5 = 1'b1;
  assign CLBLL_R_X81Y111_SLICE_X127Y111_D6 = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_T1 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_D1 = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign LIOB33_X0Y195_IOB_X0Y196_O = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign LIOB33_X0Y195_IOB_X0Y195_O = 1'b0;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B6 = CLBLM_R_X15Y114_SLICE_X20Y114_AO5;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_T1 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C5 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_T1 = 1'b1;
  assign LIOI3_X0Y85_ILOGIC_X0Y86_D = LIOB33_X0Y85_IOB_X0Y86_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_D = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C4 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C5 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLL_L_X2Y174_SLICE_X0Y174_AO5;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C6 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_D1 = CLBLM_R_X103Y103_SLICE_X163Y103_AO6;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_T1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign RIOB33_X105Y59_IOB_X1Y60_O = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign RIOB33_X105Y59_IOB_X1Y59_O = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLM_R_X93Y122_SLICE_X147Y122_CO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOB33_X0Y197_IOB_X0Y198_O = CLBLL_L_X2Y101_SLICE_X0Y101_BO6;
  assign LIOB33_X0Y197_IOB_X0Y197_O = CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_D1 = CLBLL_R_X81Y111_SLICE_X126Y111_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_R_X101Y124_SLICE_X158Y124_BO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_T1 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A4 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_D1 = CLBLM_R_X37Y111_SLICE_X56Y111_BO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1 = CLBLM_R_X15Y110_SLICE_X20Y110_DO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1 = CLBLM_R_X103Y103_SLICE_X163Y103_BO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A2 = RIOB33_X105Y153_IOB_X1Y154_I;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B4 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B5 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A3 = RIOB33_X105Y153_IOB_X1Y153_I;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A4 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C2 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C3 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C4 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A2 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A3 = RIOB33_X105Y155_IOB_X1Y156_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A4 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A5 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D6 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B2 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B3 = RIOB33_X105Y159_IOB_X1Y160_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B4 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B5 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C2 = CLBLM_R_X13Y111_SLICE_X19Y111_AO5;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C3 = CLBLM_R_X15Y111_SLICE_X21Y111_BO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C4 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C5 = RIOB33_X105Y159_IOB_X1Y160_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C6 = CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_D = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_D = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D1 = CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D2 = CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D3 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D4 = CLBLM_R_X15Y113_SLICE_X21Y113_AO5;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D5 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D6 = CLBLM_R_X15Y113_SLICE_X20Y113_AO6;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y90_D = LIOB33_X0Y89_IOB_X0Y90_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y89_D = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A1 = LIOB33_X0Y91_IOB_X0Y92_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A3 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A4 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A5 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y166_D = RIOB33_X105Y165_IOB_X1Y166_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B2 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B3 = RIOB33_X105Y157_IOB_X1Y158_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B4 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C1 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C2 = CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C3 = RIOB33_X105Y171_IOB_X1Y172_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C4 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C5 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D1 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D2 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D3 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D5 = RIOB33_X105Y157_IOB_X1Y158_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D6 = CLBLM_R_X15Y113_SLICE_X20Y113_BO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C3 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = CLBLL_L_X2Y136_SLICE_X0Y136_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = CLBLL_L_X2Y101_SLICE_X0Y101_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_D = RIOB33_X105Y157_IOB_X1Y158_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_D = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B1 = 1'b1;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_D = LIOB33_X0Y147_IOB_X0Y147_I;
  assign LIOI3_SING_X0Y99_ILOGIC_X0Y99_D = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A1 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A2 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A3 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A4 = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A6 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLM_L_X78Y125_SLICE_X121Y125_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B3 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B6 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B4 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B5 = CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_A2 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_A3 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_A5 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_A6 = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_B1 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A1 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A2 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A3 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A4 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A5 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_B2 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_B3 = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_B4 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B1 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B2 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B3 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B4 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B5 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_C1 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_C2 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C1 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C2 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C3 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C4 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C5 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_D1 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_D2 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_D3 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_D4 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_D5 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X163Y103_D6 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D1 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D2 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D3 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D4 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D5 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C5 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_A1 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_A2 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C6 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_A3 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_A4 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A2 = RIOB33_X105Y159_IOB_X1Y159_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A3 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A4 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A6 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_B1 = 1'b1;
  assign CLBLM_R_X103Y103_SLICE_X162Y103_B2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B1 = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B2 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B5 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C1 = CLBLM_R_X15Y114_SLICE_X20Y114_AO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C2 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C3 = RIOB33_X105Y159_IOB_X1Y159_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C5 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C6 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = RIOB33_X105Y161_IOB_X1Y161_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D1 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D3 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D5 = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D6 = CLBLM_R_X15Y114_SLICE_X20Y114_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = CLBLL_L_X2Y101_SLICE_X0Y101_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D6 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A1 = CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A3 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A4 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A6 = CLBLM_R_X93Y116_SLICE_X147Y116_AO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B1 = CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B3 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B4 = CLBLM_R_X93Y116_SLICE_X147Y116_AO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B5 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B6 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C6 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign RIOB33_X105Y51_IOB_X1Y52_O = CLBLM_R_X15Y99_SLICE_X20Y99_AO6;
  assign RIOB33_X105Y51_IOB_X1Y51_O = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLL_L_X2Y174_SLICE_X0Y174_AO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = CLBLM_L_X94Y122_SLICE_X148Y122_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLL_L_X2Y174_SLICE_X0Y174_AO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_D1 = CLBLM_R_X37Y111_SLICE_X56Y111_CO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLM_L_X78Y119_SLICE_X121Y119_CO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_D1 = CLBLM_L_X30Y111_SLICE_X44Y111_AO6;
  assign LIOB33_X0Y185_IOB_X0Y185_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A1 = CLBLM_R_X15Y113_SLICE_X21Y113_BO5;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A2 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A4 = CLBLM_R_X15Y111_SLICE_X21Y111_BO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A5 = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B2 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D2 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A2 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C2 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D2 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D6 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A1 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A3 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A4 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A5 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A6 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B5 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B6 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D6 = 1'b1;
  assign RIOB33_SING_X105Y50_IOB_X1Y50_O = CLBLM_R_X15Y99_SLICE_X20Y99_AO6;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_D = RIOB33_X105Y169_IOB_X1Y170_I;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_D = RIOB33_X105Y169_IOB_X1Y169_I;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B6 = 1'b1;
  assign RIOB33_X105Y53_IOB_X1Y53_O = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign RIOB33_X105Y53_IOB_X1Y54_O = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C6 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLM_L_X78Y119_SLICE_X121Y119_AO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B4 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y174_SLICE_X1Y174_D5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  assign RIOB33_SING_X105Y99_IOB_X1Y99_O = CLBLM_L_X78Y119_SLICE_X121Y119_BO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C4 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C5 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D5 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = 1'b1;
  assign RIOB33_X105Y55_IOB_X1Y56_O = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = 1'b1;
  assign RIOB33_X105Y55_IOB_X1Y55_O = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_B6 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_C3 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_C4 = 1'b1;
  assign CLBLM_R_X37Y111_SLICE_X57Y111_C6 = 1'b1;
endmodule
